
module clk_buf (
	dout,
	pad_in);	

	output	[0:0]	dout;
	input	[0:0]	pad_in;
endmodule
