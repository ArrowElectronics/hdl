
module clk2 (
	rst,
	refclk,
	outclk_0,
	outclk_1);	

	input		rst;
	input		refclk;
	output		outclk_0;
	output		outclk_1;
endmodule
