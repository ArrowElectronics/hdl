// system_bd.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module system_bd (
		output wire        hdmi_out_h_clk,                              //                        hdmi_out.h_clk
		output wire        hdmi_out_h16_hsync,                          //                                .h16_hsync
		output wire        hdmi_out_h16_vsync,                          //                                .h16_vsync
		output wire        hdmi_out_h16_data_e,                         //                                .h16_data_e
		output wire [15:0] hdmi_out_h16_data,                           //                                .h16_data
		output wire [15:0] hdmi_out_h16_es_data,                        //                                .h16_es_data
		output wire        hdmi_out_h24_hsync,                          //                                .h24_hsync
		output wire        hdmi_out_h24_vsync,                          //                                .h24_vsync
		output wire        hdmi_out_h24_data_e,                         //                                .h24_data_e
		output wire [23:0] hdmi_out_h24_data,                           //                                .h24_data
		output wire        hdmi_out_h36_hsync,                          //                                .h36_hsync
		output wire        hdmi_out_h36_vsync,                          //                                .h36_vsync
		output wire        hdmi_out_h36_data_e,                         //                                .h36_data_e
		output wire [35:0] hdmi_out_h36_data,                           //                                .h36_data
		output wire        spi_engine_execution_0_spi_out_three_wire,   //  spi_engine_execution_0_spi_out.three_wire
		output wire        spi_engine_execution_0_spi_out_sdo_t,        //                                .sdo_t
		output wire        spi_engine_execution_0_spi_out_sdo,          //                                .sdo
		input  wire        spi_engine_execution_0_spi_out_sdi,          //                                .sdi
		output wire [0:0]  spi_engine_execution_0_spi_out_cs,           //                                .cs
		output wire        spi_engine_execution_0_spi_out_sclk,         //                                .sclk
		input  wire        spi_engine_execution_0_spi_out_sdi_1,        //                                .sdi_1
		input  wire        sys_clk_clk,                                 //                         sys_clk.clk
		input  wire [31:0] sys_gpio_bd_in_port,                         //                     sys_gpio_bd.in_port
		output wire [31:0] sys_gpio_bd_out_port,                        //                                .out_port
		input  wire [31:0] sys_gpio_in_export,                          //                     sys_gpio_in.export
		output wire [31:0] sys_gpio_out_export,                         //                    sys_gpio_out.export
		output wire        sys_hps_h2f_reset_reset_n,                   //               sys_hps_h2f_reset.reset_n
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TX_CLK,     //                  sys_hps_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD0,       //                                .hps_io_emac1_inst_TXD0
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD1,       //                                .hps_io_emac1_inst_TXD1
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD2,       //                                .hps_io_emac1_inst_TXD2
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD3,       //                                .hps_io_emac1_inst_TXD3
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD0,       //                                .hps_io_emac1_inst_RXD0
		inout  wire        sys_hps_hps_io_hps_io_emac1_inst_MDIO,       //                                .hps_io_emac1_inst_MDIO
		output wire        sys_hps_hps_io_hps_io_emac1_inst_MDC,        //                                .hps_io_emac1_inst_MDC
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RX_CTL,     //                                .hps_io_emac1_inst_RX_CTL
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TX_CTL,     //                                .hps_io_emac1_inst_TX_CTL
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RX_CLK,     //                                .hps_io_emac1_inst_RX_CLK
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD1,       //                                .hps_io_emac1_inst_RXD1
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD2,       //                                .hps_io_emac1_inst_RXD2
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD3,       //                                .hps_io_emac1_inst_RXD3
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO0,         //                                .hps_io_qspi_inst_IO0
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO1,         //                                .hps_io_qspi_inst_IO1
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO2,         //                                .hps_io_qspi_inst_IO2
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO3,         //                                .hps_io_qspi_inst_IO3
		output wire        sys_hps_hps_io_hps_io_qspi_inst_SS0,         //                                .hps_io_qspi_inst_SS0
		output wire        sys_hps_hps_io_hps_io_qspi_inst_CLK,         //                                .hps_io_qspi_inst_CLK
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_CMD,         //                                .hps_io_sdio_inst_CMD
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D0,          //                                .hps_io_sdio_inst_D0
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D1,          //                                .hps_io_sdio_inst_D1
		output wire        sys_hps_hps_io_hps_io_sdio_inst_CLK,         //                                .hps_io_sdio_inst_CLK
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D2,          //                                .hps_io_sdio_inst_D2
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D3,          //                                .hps_io_sdio_inst_D3
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D0,          //                                .hps_io_usb1_inst_D0
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D1,          //                                .hps_io_usb1_inst_D1
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D2,          //                                .hps_io_usb1_inst_D2
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D3,          //                                .hps_io_usb1_inst_D3
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D4,          //                                .hps_io_usb1_inst_D4
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D5,          //                                .hps_io_usb1_inst_D5
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D6,          //                                .hps_io_usb1_inst_D6
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D7,          //                                .hps_io_usb1_inst_D7
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_CLK,         //                                .hps_io_usb1_inst_CLK
		output wire        sys_hps_hps_io_hps_io_usb1_inst_STP,         //                                .hps_io_usb1_inst_STP
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_DIR,         //                                .hps_io_usb1_inst_DIR
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_NXT,         //                                .hps_io_usb1_inst_NXT
		input  wire        sys_hps_hps_io_hps_io_uart0_inst_RX,         //                                .hps_io_uart0_inst_RX
		output wire        sys_hps_hps_io_hps_io_uart0_inst_TX,         //                                .hps_io_uart0_inst_TX
		inout  wire        sys_hps_hps_io_hps_io_i2c0_inst_SDA,         //                                .hps_io_i2c0_inst_SDA
		inout  wire        sys_hps_hps_io_hps_io_i2c0_inst_SCL,         //                                .hps_io_i2c0_inst_SCL
		inout  wire        sys_hps_hps_io_hps_io_i2c1_inst_SDA,         //                                .hps_io_i2c1_inst_SDA
		inout  wire        sys_hps_hps_io_hps_io_i2c1_inst_SCL,         //                                .hps_io_i2c1_inst_SCL
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO00,      //                                .hps_io_gpio_inst_GPIO00
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO09,      //                                .hps_io_gpio_inst_GPIO09
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO35,      //                                .hps_io_gpio_inst_GPIO35
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO40,      //                                .hps_io_gpio_inst_GPIO40
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO41,      //                                .hps_io_gpio_inst_GPIO41
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO42,      //                                .hps_io_gpio_inst_GPIO42
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO43,      //                                .hps_io_gpio_inst_GPIO43
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO44,      //                                .hps_io_gpio_inst_GPIO44
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO48,      //                                .hps_io_gpio_inst_GPIO48
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO53,      //                                .hps_io_gpio_inst_GPIO53
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO54,      //                                .hps_io_gpio_inst_GPIO54
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO55,      //                                .hps_io_gpio_inst_GPIO55
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO56,      //                                .hps_io_gpio_inst_GPIO56
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO57,      //                                .hps_io_gpio_inst_GPIO57
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO58,      //                                .hps_io_gpio_inst_GPIO58
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO59,      //                                .hps_io_gpio_inst_GPIO59
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO61,      //                                .hps_io_gpio_inst_GPIO61
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO65,      //                                .hps_io_gpio_inst_GPIO65
		output wire [15:0] sys_hps_memory_mem_a,                        //                  sys_hps_memory.mem_a
		output wire [2:0]  sys_hps_memory_mem_ba,                       //                                .mem_ba
		output wire        sys_hps_memory_mem_ck,                       //                                .mem_ck
		output wire        sys_hps_memory_mem_ck_n,                     //                                .mem_ck_n
		output wire        sys_hps_memory_mem_cke,                      //                                .mem_cke
		output wire        sys_hps_memory_mem_cs_n,                     //                                .mem_cs_n
		output wire        sys_hps_memory_mem_ras_n,                    //                                .mem_ras_n
		output wire        sys_hps_memory_mem_cas_n,                    //                                .mem_cas_n
		output wire        sys_hps_memory_mem_we_n,                     //                                .mem_we_n
		output wire        sys_hps_memory_mem_reset_n,                  //                                .mem_reset_n
		inout  wire [31:0] sys_hps_memory_mem_dq,                       //                                .mem_dq
		inout  wire [3:0]  sys_hps_memory_mem_dqs,                      //                                .mem_dqs
		inout  wire [3:0]  sys_hps_memory_mem_dqs_n,                    //                                .mem_dqs_n
		output wire        sys_hps_memory_mem_odt,                      //                                .mem_odt
		output wire [3:0]  sys_hps_memory_mem_dm,                       //                                .mem_dm
		input  wire        sys_hps_memory_oct_rzqin,                    //                                .oct_rzqin
		input  wire        sys_rst_reset_n,                             //                         sys_rst.reset_n
		input  wire        trigger_gen_0_load_config_load_config,       //       trigger_gen_0_load_config.load_config
		input  wire [31:0] trigger_gen_0_pulse_period_pulse_period,     //      trigger_gen_0_pulse_period.pulse_period
		input  wire [31:0] trigger_gen_0_pulse_width_pulse_width,       //       trigger_gen_0_pulse_width.pulse_width
		input  wire        upscale_converter_0_dfmt_enable_dfmt_enable, // upscale_converter_0_dfmt_enable.dfmt_enable
		input  wire        upscale_converter_0_dfmt_se_dfmt_se,         //     upscale_converter_0_dfmt_se.dfmt_se
		input  wire        upscale_converter_0_dfmt_type_dfmt_type      //   upscale_converter_0_dfmt_type.dfmt_type
	);

	wire         upscale_converter_0_m_axis_tvalid;                       // upscale_converter_0:m_axis_valid -> spi_dmac_0:s_axis_valid
	wire         upscale_converter_0_m_axis_tready;                       // spi_dmac_0:s_axis_ready -> upscale_converter_0:m_axis_ready
	wire  [63:0] upscale_converter_0_m_axis_tdata;                        // upscale_converter_0:m_axis_data -> spi_dmac_0:s_axis_data
	wire         hdmi_dmac_0_m_axis_tvalid;                               // hdmi_dmac_0:m_axis_valid -> axi_hdmi_tx_0:vdma_valid
	wire         hdmi_dmac_0_m_axis_tready;                               // axi_hdmi_tx_0:vdma_ready -> hdmi_dmac_0:m_axis_ready
	wire         hdmi_dmac_0_m_axis_tlast;                                // hdmi_dmac_0:m_axis_last -> axi_hdmi_tx_0:vdma_end_of_frame
	wire  [63:0] hdmi_dmac_0_m_axis_tdata;                                // hdmi_dmac_0:m_axis_data -> axi_hdmi_tx_0:vdma_data
	wire         sys_hps_h2f_user1_clock_clk;                             // sys_hps:h2f_user1_clk -> [axi_hdmi_tx_0:s_axi_aclk, axi_hdmi_tx_0:vdma_clk, axi_spi_engine_0:s_axi_aclk, hdmi_dmac_0:m_axis_aclk, hdmi_dmac_0:m_src_axi_aclk, hdmi_dmac_0:s_axi_aclk, hdmi_pll:refclk, mm_interconnect_0:sys_hps_h2f_user1_clock_clk, mm_interconnect_1:sys_hps_h2f_user1_clock_clk, mm_interconnect_2:sys_hps_h2f_user1_clock_clk, rst_controller:clk, rst_controller_001:clk, spi_dmac_0:m_dest_axi_aclk, spi_dmac_0:s_axi_aclk, spi_engine_pll:refclk, sys_gpio_bd:clk, sys_gpio_in:clk, sys_gpio_out:clk, sys_hps:f2h_axi_clk, sys_hps:f2h_sdram0_clk, sys_hps:f2h_sdram1_clk, sys_hps:f2h_sdram2_clk, sys_hps:h2f_axi_clk, sys_hps:h2f_lw_axi_clk, sys_id:clock]
	wire         spi_engine_pll_outclk0_clk;                              // spi_engine_pll:outclk_0 -> [axi_spi_engine_0:spi_clk, spi_dmac_0:s_axis_aclk, spi_engine_execution_0:clk, spi_engine_interconnect_0:clk, spi_engine_offload_0:ctrl_clk, spi_engine_offload_0:spi_clk, trigger_gen_0:clk, upscale_converter_0:clk]
	wire         hdmi_pll_outclk0_clk;                                    // hdmi_pll:outclk_0 -> axi_hdmi_tx_0:hdmi_clk
	wire         spi_engine_execution_0_ctrl_sync_valid;                  // spi_engine_execution_0:sync_valid -> spi_engine_interconnect_0:m_sync_valid
	wire  [17:0] spi_engine_interconnect_0_m_ctrl_sdo_data;               // spi_engine_interconnect_0:m_sdo_data -> spi_engine_execution_0:sdo_data
	wire         spi_engine_interconnect_0_m_ctrl_sdi_data_ready;         // spi_engine_interconnect_0:m_sdi_ready -> spi_engine_execution_0:sdi_data_ready
	wire         spi_engine_execution_0_ctrl_sdo_data_ready;              // spi_engine_execution_0:sdo_data_ready -> spi_engine_interconnect_0:m_sdo_ready
	wire         spi_engine_execution_0_ctrl_cmd_ready;                   // spi_engine_execution_0:cmd_ready -> spi_engine_interconnect_0:m_cmd_ready
	wire         spi_engine_interconnect_0_m_ctrl_cmd_valid;              // spi_engine_interconnect_0:m_cmd_valid -> spi_engine_execution_0:cmd_valid
	wire         spi_engine_interconnect_0_m_ctrl_sdo_data_valid;         // spi_engine_interconnect_0:m_sdo_valid -> spi_engine_execution_0:sdo_data_valid
	wire         spi_engine_execution_0_ctrl_sdi_data_valid;              // spi_engine_execution_0:sdi_data_valid -> spi_engine_interconnect_0:m_sdi_valid
	wire  [15:0] spi_engine_interconnect_0_m_ctrl_cmd;                    // spi_engine_interconnect_0:m_cmd_data -> spi_engine_execution_0:cmd
	wire  [35:0] spi_engine_execution_0_ctrl_sdi_data;                    // spi_engine_execution_0:sdi_data -> spi_engine_interconnect_0:m_sdi_data
	wire   [7:0] spi_engine_execution_0_ctrl_sync;                        // spi_engine_execution_0:sync -> spi_engine_interconnect_0:m_sync
	wire         spi_engine_interconnect_0_m_ctrl_sync_ready;             // spi_engine_interconnect_0:m_sync_ready -> spi_engine_execution_0:sync_ready
	wire         spi_engine_offload_0_offload_sdi_valid;                  // spi_engine_offload_0:offload_sdi_valid -> upscale_converter_0:s_axis_valid
	wire  [35:0] spi_engine_offload_0_offload_sdi_data;                   // spi_engine_offload_0:offload_sdi_data -> upscale_converter_0:s_axis_data
	wire         upscale_converter_0_s_axis_ready;                        // upscale_converter_0:s_axis_ready -> spi_engine_offload_0:offload_sdi_ready
	wire         trigger_gen_0_pulse_pulse;                               // trigger_gen_0:pulse -> spi_engine_offload_0:trigger
	wire         spi_engine_interconnect_0_s0_ctrl_sync_valid;            // spi_engine_interconnect_0:s0_sync_valid -> spi_engine_offload_0:sync_valid
	wire  [17:0] spi_engine_offload_0_spi_engine_ctrl_sdo_data;           // spi_engine_offload_0:sdo_data -> spi_engine_interconnect_0:s0_sdo_data
	wire         spi_engine_interconnect_0_s0_ctrl_cmd_ready;             // spi_engine_interconnect_0:s0_cmd_ready -> spi_engine_offload_0:cmd_ready
	wire  [15:0] spi_engine_offload_0_spi_engine_ctrl_cmd_data;           // spi_engine_offload_0:cmd -> spi_engine_interconnect_0:s0_cmd_data
	wire         spi_engine_offload_0_spi_engine_ctrl_cmd_valid;          // spi_engine_offload_0:cmd_valid -> spi_engine_interconnect_0:s0_cmd_valid
	wire         spi_engine_interconnect_0_s0_ctrl_sdo_ready;             // spi_engine_interconnect_0:s0_sdo_ready -> spi_engine_offload_0:sdo_data_ready
	wire         spi_engine_offload_0_spi_engine_ctrl_sdo_valid;          // spi_engine_offload_0:sdo_data_valid -> spi_engine_interconnect_0:s0_sdo_valid
	wire   [7:0] spi_engine_interconnect_0_s0_ctrl_sync_data;             // spi_engine_interconnect_0:s0_sync -> spi_engine_offload_0:sync_data
	wire  [35:0] spi_engine_interconnect_0_s0_ctrl_sdi_data;              // spi_engine_interconnect_0:s0_sdi_data -> spi_engine_offload_0:sdi_data
	wire         spi_engine_offload_0_spi_engine_ctrl_sync_ready;         // spi_engine_offload_0:sync_ready -> spi_engine_interconnect_0:s0_sync_ready
	wire         spi_engine_offload_0_spi_engine_ctrl_sdi_ready;          // spi_engine_offload_0:sdi_data_ready -> spi_engine_interconnect_0:s0_sdi_ready
	wire         spi_engine_interconnect_0_s0_ctrl_sdi_valid;             // spi_engine_interconnect_0:s0_sdi_valid -> spi_engine_offload_0:sdi_data_valid
	wire         spi_engine_interconnect_0_s1_ctrl_sync_valid;            // spi_engine_interconnect_0:s1_sync_valid -> axi_spi_engine_0:sync_valid
	wire  [17:0] axi_spi_engine_0_spi_engine_ctrl_sdo_data;               // axi_spi_engine_0:sdo_data -> spi_engine_interconnect_0:s1_sdo_data
	wire         spi_engine_interconnect_0_s1_ctrl_cmd_ready;             // spi_engine_interconnect_0:s1_cmd_ready -> axi_spi_engine_0:cmd_ready
	wire  [15:0] axi_spi_engine_0_spi_engine_ctrl_cmd_data;               // axi_spi_engine_0:cmd_data -> spi_engine_interconnect_0:s1_cmd_data
	wire         axi_spi_engine_0_spi_engine_ctrl_cmd_valid;              // axi_spi_engine_0:cmd_valid -> spi_engine_interconnect_0:s1_cmd_valid
	wire         spi_engine_interconnect_0_s1_ctrl_sdo_ready;             // spi_engine_interconnect_0:s1_sdo_ready -> axi_spi_engine_0:sdo_data_ready
	wire         axi_spi_engine_0_spi_engine_ctrl_sdo_valid;              // axi_spi_engine_0:sdo_data_valid -> spi_engine_interconnect_0:s1_sdo_valid
	wire   [7:0] spi_engine_interconnect_0_s1_ctrl_sync_data;             // spi_engine_interconnect_0:s1_sync -> axi_spi_engine_0:sync_data
	wire  [35:0] spi_engine_interconnect_0_s1_ctrl_sdi_data;              // spi_engine_interconnect_0:s1_sdi_data -> axi_spi_engine_0:sdi_data
	wire         axi_spi_engine_0_spi_engine_ctrl_sync_ready;             // axi_spi_engine_0:sync_ready -> spi_engine_interconnect_0:s1_sync_ready
	wire         axi_spi_engine_0_spi_engine_ctrl_sdi_ready;              // axi_spi_engine_0:sdi_data_ready -> spi_engine_interconnect_0:s1_sdi_ready
	wire         spi_engine_interconnect_0_s1_ctrl_sdi_valid;             // spi_engine_interconnect_0:s1_sdi_valid -> axi_spi_engine_0:sdi_data_valid
	wire  [15:0] axi_spi_engine_0_spi_engine_offload_ctrl0_cmd_wr_data;   // axi_spi_engine_0:offload0_cmd_wr_data -> spi_engine_offload_0:ctrl_cmd_wr_data
	wire  [17:0] axi_spi_engine_0_spi_engine_offload_ctrl0_sdo_wr_data;   // axi_spi_engine_0:offload0_sdo_wr_data -> spi_engine_offload_0:ctrl_sdo_wr_data
	wire         axi_spi_engine_0_spi_engine_offload_ctrl0_enable;        // axi_spi_engine_0:offload0_enable -> spi_engine_offload_0:ctrl_enable
	wire         axi_spi_engine_0_spi_engine_offload_ctrl0_sdo_wr_en;     // axi_spi_engine_0:offload0_sdo_wr_en -> spi_engine_offload_0:ctrl_sdo_wr_en
	wire         axi_spi_engine_0_spi_engine_offload_ctrl0_reset;         // axi_spi_engine_0:offload0_mem_reset -> spi_engine_offload_0:ctrl_mem_reset
	wire         axi_spi_engine_0_spi_engine_offload_ctrl0_cmd_wr_en;     // axi_spi_engine_0:offload0_cmd_wr_en -> spi_engine_offload_0:ctrl_cmd_wr_en
	wire         spi_engine_offload_0_spi_engine_offload_ctrl_enabled;    // spi_engine_offload_0:ctrl_enabled -> axi_spi_engine_0:offload0_enabled
	wire         axi_spi_engine_0_spi_resetn_reset;                       // axi_spi_engine_0:spi_resetn -> [spi_engine_execution_0:resetn, spi_engine_interconnect_0:resetn, spi_engine_offload_0:spi_resetn, trigger_gen_0:rstn, upscale_converter_0:resetn]
	wire   [1:0] sys_hps_h2f_lw_axi_master_awburst;                       // sys_hps:h2f_lw_AWBURST -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awburst
	wire   [3:0] sys_hps_h2f_lw_axi_master_arlen;                         // sys_hps:h2f_lw_ARLEN -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arlen
	wire   [3:0] sys_hps_h2f_lw_axi_master_wstrb;                         // sys_hps:h2f_lw_WSTRB -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wstrb
	wire         sys_hps_h2f_lw_axi_master_wready;                        // mm_interconnect_0:sys_hps_h2f_lw_axi_master_wready -> sys_hps:h2f_lw_WREADY
	wire  [11:0] sys_hps_h2f_lw_axi_master_rid;                           // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rid -> sys_hps:h2f_lw_RID
	wire         sys_hps_h2f_lw_axi_master_rready;                        // sys_hps:h2f_lw_RREADY -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_rready
	wire   [3:0] sys_hps_h2f_lw_axi_master_awlen;                         // sys_hps:h2f_lw_AWLEN -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awlen
	wire  [11:0] sys_hps_h2f_lw_axi_master_wid;                           // sys_hps:h2f_lw_WID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wid
	wire   [3:0] sys_hps_h2f_lw_axi_master_arcache;                       // sys_hps:h2f_lw_ARCACHE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arcache
	wire         sys_hps_h2f_lw_axi_master_wvalid;                        // sys_hps:h2f_lw_WVALID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wvalid
	wire  [20:0] sys_hps_h2f_lw_axi_master_araddr;                        // sys_hps:h2f_lw_ARADDR -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_araddr
	wire   [2:0] sys_hps_h2f_lw_axi_master_arprot;                        // sys_hps:h2f_lw_ARPROT -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arprot
	wire   [2:0] sys_hps_h2f_lw_axi_master_awprot;                        // sys_hps:h2f_lw_AWPROT -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awprot
	wire  [31:0] sys_hps_h2f_lw_axi_master_wdata;                         // sys_hps:h2f_lw_WDATA -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wdata
	wire         sys_hps_h2f_lw_axi_master_arvalid;                       // sys_hps:h2f_lw_ARVALID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arvalid
	wire   [3:0] sys_hps_h2f_lw_axi_master_awcache;                       // sys_hps:h2f_lw_AWCACHE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awcache
	wire  [11:0] sys_hps_h2f_lw_axi_master_arid;                          // sys_hps:h2f_lw_ARID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arid
	wire   [1:0] sys_hps_h2f_lw_axi_master_arlock;                        // sys_hps:h2f_lw_ARLOCK -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arlock
	wire   [1:0] sys_hps_h2f_lw_axi_master_awlock;                        // sys_hps:h2f_lw_AWLOCK -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awlock
	wire  [20:0] sys_hps_h2f_lw_axi_master_awaddr;                        // sys_hps:h2f_lw_AWADDR -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awaddr
	wire   [1:0] sys_hps_h2f_lw_axi_master_bresp;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_bresp -> sys_hps:h2f_lw_BRESP
	wire         sys_hps_h2f_lw_axi_master_arready;                       // mm_interconnect_0:sys_hps_h2f_lw_axi_master_arready -> sys_hps:h2f_lw_ARREADY
	wire  [31:0] sys_hps_h2f_lw_axi_master_rdata;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rdata -> sys_hps:h2f_lw_RDATA
	wire         sys_hps_h2f_lw_axi_master_awready;                       // mm_interconnect_0:sys_hps_h2f_lw_axi_master_awready -> sys_hps:h2f_lw_AWREADY
	wire   [1:0] sys_hps_h2f_lw_axi_master_arburst;                       // sys_hps:h2f_lw_ARBURST -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arburst
	wire   [2:0] sys_hps_h2f_lw_axi_master_arsize;                        // sys_hps:h2f_lw_ARSIZE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arsize
	wire         sys_hps_h2f_lw_axi_master_bready;                        // sys_hps:h2f_lw_BREADY -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_bready
	wire         sys_hps_h2f_lw_axi_master_rlast;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rlast -> sys_hps:h2f_lw_RLAST
	wire         sys_hps_h2f_lw_axi_master_wlast;                         // sys_hps:h2f_lw_WLAST -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wlast
	wire   [1:0] sys_hps_h2f_lw_axi_master_rresp;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rresp -> sys_hps:h2f_lw_RRESP
	wire  [11:0] sys_hps_h2f_lw_axi_master_awid;                          // sys_hps:h2f_lw_AWID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awid
	wire  [11:0] sys_hps_h2f_lw_axi_master_bid;                           // mm_interconnect_0:sys_hps_h2f_lw_axi_master_bid -> sys_hps:h2f_lw_BID
	wire         sys_hps_h2f_lw_axi_master_bvalid;                        // mm_interconnect_0:sys_hps_h2f_lw_axi_master_bvalid -> sys_hps:h2f_lw_BVALID
	wire   [2:0] sys_hps_h2f_lw_axi_master_awsize;                        // sys_hps:h2f_lw_AWSIZE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awsize
	wire         sys_hps_h2f_lw_axi_master_awvalid;                       // sys_hps:h2f_lw_AWVALID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awvalid
	wire         sys_hps_h2f_lw_axi_master_rvalid;                        // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rvalid -> sys_hps:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;         // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;          // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire         mm_interconnect_0_sys_gpio_bd_s1_chipselect;             // mm_interconnect_0:sys_gpio_bd_s1_chipselect -> sys_gpio_bd:chipselect
	wire  [31:0] mm_interconnect_0_sys_gpio_bd_s1_readdata;               // sys_gpio_bd:readdata -> mm_interconnect_0:sys_gpio_bd_s1_readdata
	wire   [1:0] mm_interconnect_0_sys_gpio_bd_s1_address;                // mm_interconnect_0:sys_gpio_bd_s1_address -> sys_gpio_bd:address
	wire         mm_interconnect_0_sys_gpio_bd_s1_write;                  // mm_interconnect_0:sys_gpio_bd_s1_write -> sys_gpio_bd:write_n
	wire  [31:0] mm_interconnect_0_sys_gpio_bd_s1_writedata;              // mm_interconnect_0:sys_gpio_bd_s1_writedata -> sys_gpio_bd:writedata
	wire         mm_interconnect_0_sys_gpio_in_s1_chipselect;             // mm_interconnect_0:sys_gpio_in_s1_chipselect -> sys_gpio_in:chipselect
	wire  [31:0] mm_interconnect_0_sys_gpio_in_s1_readdata;               // sys_gpio_in:readdata -> mm_interconnect_0:sys_gpio_in_s1_readdata
	wire   [1:0] mm_interconnect_0_sys_gpio_in_s1_address;                // mm_interconnect_0:sys_gpio_in_s1_address -> sys_gpio_in:address
	wire         mm_interconnect_0_sys_gpio_in_s1_write;                  // mm_interconnect_0:sys_gpio_in_s1_write -> sys_gpio_in:write_n
	wire  [31:0] mm_interconnect_0_sys_gpio_in_s1_writedata;              // mm_interconnect_0:sys_gpio_in_s1_writedata -> sys_gpio_in:writedata
	wire         mm_interconnect_0_sys_gpio_out_s1_chipselect;            // mm_interconnect_0:sys_gpio_out_s1_chipselect -> sys_gpio_out:chipselect
	wire  [31:0] mm_interconnect_0_sys_gpio_out_s1_readdata;              // sys_gpio_out:readdata -> mm_interconnect_0:sys_gpio_out_s1_readdata
	wire   [1:0] mm_interconnect_0_sys_gpio_out_s1_address;               // mm_interconnect_0:sys_gpio_out_s1_address -> sys_gpio_out:address
	wire         mm_interconnect_0_sys_gpio_out_s1_write;                 // mm_interconnect_0:sys_gpio_out_s1_write -> sys_gpio_out:write_n
	wire  [31:0] mm_interconnect_0_sys_gpio_out_s1_writedata;             // mm_interconnect_0:sys_gpio_out_s1_writedata -> sys_gpio_out:writedata
	wire  [10:0] mm_interconnect_0_hdmi_dmac_0_s_axi_awaddr;              // mm_interconnect_0:hdmi_dmac_0_s_axi_awaddr -> hdmi_dmac_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_hdmi_dmac_0_s_axi_bresp;               // hdmi_dmac_0:s_axi_bresp -> mm_interconnect_0:hdmi_dmac_0_s_axi_bresp
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_arready;             // hdmi_dmac_0:s_axi_arready -> mm_interconnect_0:hdmi_dmac_0_s_axi_arready
	wire  [31:0] mm_interconnect_0_hdmi_dmac_0_s_axi_rdata;               // hdmi_dmac_0:s_axi_rdata -> mm_interconnect_0:hdmi_dmac_0_s_axi_rdata
	wire   [3:0] mm_interconnect_0_hdmi_dmac_0_s_axi_wstrb;               // mm_interconnect_0:hdmi_dmac_0_s_axi_wstrb -> hdmi_dmac_0:s_axi_wstrb
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_wready;              // hdmi_dmac_0:s_axi_wready -> mm_interconnect_0:hdmi_dmac_0_s_axi_wready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_awready;             // hdmi_dmac_0:s_axi_awready -> mm_interconnect_0:hdmi_dmac_0_s_axi_awready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_rready;              // mm_interconnect_0:hdmi_dmac_0_s_axi_rready -> hdmi_dmac_0:s_axi_rready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_bready;              // mm_interconnect_0:hdmi_dmac_0_s_axi_bready -> hdmi_dmac_0:s_axi_bready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_wvalid;              // mm_interconnect_0:hdmi_dmac_0_s_axi_wvalid -> hdmi_dmac_0:s_axi_wvalid
	wire  [10:0] mm_interconnect_0_hdmi_dmac_0_s_axi_araddr;              // mm_interconnect_0:hdmi_dmac_0_s_axi_araddr -> hdmi_dmac_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_hdmi_dmac_0_s_axi_arprot;              // mm_interconnect_0:hdmi_dmac_0_s_axi_arprot -> hdmi_dmac_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_hdmi_dmac_0_s_axi_rresp;               // hdmi_dmac_0:s_axi_rresp -> mm_interconnect_0:hdmi_dmac_0_s_axi_rresp
	wire   [2:0] mm_interconnect_0_hdmi_dmac_0_s_axi_awprot;              // mm_interconnect_0:hdmi_dmac_0_s_axi_awprot -> hdmi_dmac_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_hdmi_dmac_0_s_axi_wdata;               // mm_interconnect_0:hdmi_dmac_0_s_axi_wdata -> hdmi_dmac_0:s_axi_wdata
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_arvalid;             // mm_interconnect_0:hdmi_dmac_0_s_axi_arvalid -> hdmi_dmac_0:s_axi_arvalid
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_bvalid;              // hdmi_dmac_0:s_axi_bvalid -> mm_interconnect_0:hdmi_dmac_0_s_axi_bvalid
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_awvalid;             // mm_interconnect_0:hdmi_dmac_0_s_axi_awvalid -> hdmi_dmac_0:s_axi_awvalid
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_rvalid;              // hdmi_dmac_0:s_axi_rvalid -> mm_interconnect_0:hdmi_dmac_0_s_axi_rvalid
	wire  [15:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_awaddr;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_awaddr -> axi_hdmi_tx_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_bresp;             // axi_hdmi_tx_0:s_axi_bresp -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_bresp
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_arready;           // axi_hdmi_tx_0:s_axi_arready -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_arready
	wire  [31:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_rdata;             // axi_hdmi_tx_0:s_axi_rdata -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_rdata
	wire   [3:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_wstrb;             // mm_interconnect_0:axi_hdmi_tx_0_s_axi_wstrb -> axi_hdmi_tx_0:s_axi_wstrb
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_wready;            // axi_hdmi_tx_0:s_axi_wready -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_wready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_awready;           // axi_hdmi_tx_0:s_axi_awready -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_awready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_rready;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_rready -> axi_hdmi_tx_0:s_axi_rready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_bready;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_bready -> axi_hdmi_tx_0:s_axi_bready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_wvalid;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_wvalid -> axi_hdmi_tx_0:s_axi_wvalid
	wire  [15:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_araddr;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_araddr -> axi_hdmi_tx_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_arprot;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_arprot -> axi_hdmi_tx_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_rresp;             // axi_hdmi_tx_0:s_axi_rresp -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_rresp
	wire   [2:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_awprot;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_awprot -> axi_hdmi_tx_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_wdata;             // mm_interconnect_0:axi_hdmi_tx_0_s_axi_wdata -> axi_hdmi_tx_0:s_axi_wdata
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_arvalid;           // mm_interconnect_0:axi_hdmi_tx_0_s_axi_arvalid -> axi_hdmi_tx_0:s_axi_arvalid
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_bvalid;            // axi_hdmi_tx_0:s_axi_bvalid -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_bvalid
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_awvalid;           // mm_interconnect_0:axi_hdmi_tx_0_s_axi_awvalid -> axi_hdmi_tx_0:s_axi_awvalid
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_rvalid;            // axi_hdmi_tx_0:s_axi_rvalid -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_rvalid
	wire  [15:0] mm_interconnect_0_axi_spi_engine_0_s_axi_awaddr;         // mm_interconnect_0:axi_spi_engine_0_s_axi_awaddr -> axi_spi_engine_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_axi_spi_engine_0_s_axi_bresp;          // axi_spi_engine_0:s_axi_bresp -> mm_interconnect_0:axi_spi_engine_0_s_axi_bresp
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_arready;        // axi_spi_engine_0:s_axi_arready -> mm_interconnect_0:axi_spi_engine_0_s_axi_arready
	wire  [31:0] mm_interconnect_0_axi_spi_engine_0_s_axi_rdata;          // axi_spi_engine_0:s_axi_rdata -> mm_interconnect_0:axi_spi_engine_0_s_axi_rdata
	wire   [3:0] mm_interconnect_0_axi_spi_engine_0_s_axi_wstrb;          // mm_interconnect_0:axi_spi_engine_0_s_axi_wstrb -> axi_spi_engine_0:s_axi_wstrb
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_wready;         // axi_spi_engine_0:s_axi_wready -> mm_interconnect_0:axi_spi_engine_0_s_axi_wready
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_awready;        // axi_spi_engine_0:s_axi_awready -> mm_interconnect_0:axi_spi_engine_0_s_axi_awready
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_rready;         // mm_interconnect_0:axi_spi_engine_0_s_axi_rready -> axi_spi_engine_0:s_axi_rready
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_bready;         // mm_interconnect_0:axi_spi_engine_0_s_axi_bready -> axi_spi_engine_0:s_axi_bready
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_wvalid;         // mm_interconnect_0:axi_spi_engine_0_s_axi_wvalid -> axi_spi_engine_0:s_axi_wvalid
	wire  [15:0] mm_interconnect_0_axi_spi_engine_0_s_axi_araddr;         // mm_interconnect_0:axi_spi_engine_0_s_axi_araddr -> axi_spi_engine_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_axi_spi_engine_0_s_axi_arprot;         // mm_interconnect_0:axi_spi_engine_0_s_axi_arprot -> axi_spi_engine_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_axi_spi_engine_0_s_axi_rresp;          // axi_spi_engine_0:s_axi_rresp -> mm_interconnect_0:axi_spi_engine_0_s_axi_rresp
	wire   [2:0] mm_interconnect_0_axi_spi_engine_0_s_axi_awprot;         // mm_interconnect_0:axi_spi_engine_0_s_axi_awprot -> axi_spi_engine_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_axi_spi_engine_0_s_axi_wdata;          // mm_interconnect_0:axi_spi_engine_0_s_axi_wdata -> axi_spi_engine_0:s_axi_wdata
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_arvalid;        // mm_interconnect_0:axi_spi_engine_0_s_axi_arvalid -> axi_spi_engine_0:s_axi_arvalid
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_bvalid;         // axi_spi_engine_0:s_axi_bvalid -> mm_interconnect_0:axi_spi_engine_0_s_axi_bvalid
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_awvalid;        // mm_interconnect_0:axi_spi_engine_0_s_axi_awvalid -> axi_spi_engine_0:s_axi_awvalid
	wire         mm_interconnect_0_axi_spi_engine_0_s_axi_rvalid;         // axi_spi_engine_0:s_axi_rvalid -> mm_interconnect_0:axi_spi_engine_0_s_axi_rvalid
	wire  [10:0] mm_interconnect_0_spi_dmac_0_s_axi_awaddr;               // mm_interconnect_0:spi_dmac_0_s_axi_awaddr -> spi_dmac_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_spi_dmac_0_s_axi_bresp;                // spi_dmac_0:s_axi_bresp -> mm_interconnect_0:spi_dmac_0_s_axi_bresp
	wire         mm_interconnect_0_spi_dmac_0_s_axi_arready;              // spi_dmac_0:s_axi_arready -> mm_interconnect_0:spi_dmac_0_s_axi_arready
	wire  [31:0] mm_interconnect_0_spi_dmac_0_s_axi_rdata;                // spi_dmac_0:s_axi_rdata -> mm_interconnect_0:spi_dmac_0_s_axi_rdata
	wire   [3:0] mm_interconnect_0_spi_dmac_0_s_axi_wstrb;                // mm_interconnect_0:spi_dmac_0_s_axi_wstrb -> spi_dmac_0:s_axi_wstrb
	wire         mm_interconnect_0_spi_dmac_0_s_axi_wready;               // spi_dmac_0:s_axi_wready -> mm_interconnect_0:spi_dmac_0_s_axi_wready
	wire         mm_interconnect_0_spi_dmac_0_s_axi_awready;              // spi_dmac_0:s_axi_awready -> mm_interconnect_0:spi_dmac_0_s_axi_awready
	wire         mm_interconnect_0_spi_dmac_0_s_axi_rready;               // mm_interconnect_0:spi_dmac_0_s_axi_rready -> spi_dmac_0:s_axi_rready
	wire         mm_interconnect_0_spi_dmac_0_s_axi_bready;               // mm_interconnect_0:spi_dmac_0_s_axi_bready -> spi_dmac_0:s_axi_bready
	wire         mm_interconnect_0_spi_dmac_0_s_axi_wvalid;               // mm_interconnect_0:spi_dmac_0_s_axi_wvalid -> spi_dmac_0:s_axi_wvalid
	wire  [10:0] mm_interconnect_0_spi_dmac_0_s_axi_araddr;               // mm_interconnect_0:spi_dmac_0_s_axi_araddr -> spi_dmac_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_spi_dmac_0_s_axi_arprot;               // mm_interconnect_0:spi_dmac_0_s_axi_arprot -> spi_dmac_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_spi_dmac_0_s_axi_rresp;                // spi_dmac_0:s_axi_rresp -> mm_interconnect_0:spi_dmac_0_s_axi_rresp
	wire   [2:0] mm_interconnect_0_spi_dmac_0_s_axi_awprot;               // mm_interconnect_0:spi_dmac_0_s_axi_awprot -> spi_dmac_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_spi_dmac_0_s_axi_wdata;                // mm_interconnect_0:spi_dmac_0_s_axi_wdata -> spi_dmac_0:s_axi_wdata
	wire         mm_interconnect_0_spi_dmac_0_s_axi_arvalid;              // mm_interconnect_0:spi_dmac_0_s_axi_arvalid -> spi_dmac_0:s_axi_arvalid
	wire         mm_interconnect_0_spi_dmac_0_s_axi_bvalid;               // spi_dmac_0:s_axi_bvalid -> mm_interconnect_0:spi_dmac_0_s_axi_bvalid
	wire         mm_interconnect_0_spi_dmac_0_s_axi_awvalid;              // mm_interconnect_0:spi_dmac_0_s_axi_awvalid -> spi_dmac_0:s_axi_awvalid
	wire         mm_interconnect_0_spi_dmac_0_s_axi_rvalid;               // spi_dmac_0:s_axi_rvalid -> mm_interconnect_0:spi_dmac_0_s_axi_rvalid
	wire   [1:0] spi_dmac_0_m_dest_axi_awburst;                           // spi_dmac_0:m_dest_axi_awburst -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awburst
	wire   [3:0] spi_dmac_0_m_dest_axi_arlen;                             // spi_dmac_0:m_dest_axi_arlen -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arlen
	wire   [7:0] spi_dmac_0_m_dest_axi_wstrb;                             // spi_dmac_0:m_dest_axi_wstrb -> mm_interconnect_1:spi_dmac_0_m_dest_axi_wstrb
	wire         spi_dmac_0_m_dest_axi_wready;                            // mm_interconnect_1:spi_dmac_0_m_dest_axi_wready -> spi_dmac_0:m_dest_axi_wready
	wire         spi_dmac_0_m_dest_axi_rid;                               // mm_interconnect_1:spi_dmac_0_m_dest_axi_rid -> spi_dmac_0:m_dest_axi_rid
	wire         spi_dmac_0_m_dest_axi_rready;                            // spi_dmac_0:m_dest_axi_rready -> mm_interconnect_1:spi_dmac_0_m_dest_axi_rready
	wire   [3:0] spi_dmac_0_m_dest_axi_awlen;                             // spi_dmac_0:m_dest_axi_awlen -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awlen
	wire         spi_dmac_0_m_dest_axi_wid;                               // spi_dmac_0:m_dest_axi_wid -> mm_interconnect_1:spi_dmac_0_m_dest_axi_wid
	wire   [3:0] spi_dmac_0_m_dest_axi_arcache;                           // spi_dmac_0:m_dest_axi_arcache -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arcache
	wire         spi_dmac_0_m_dest_axi_wvalid;                            // spi_dmac_0:m_dest_axi_wvalid -> mm_interconnect_1:spi_dmac_0_m_dest_axi_wvalid
	wire  [31:0] spi_dmac_0_m_dest_axi_araddr;                            // spi_dmac_0:m_dest_axi_araddr -> mm_interconnect_1:spi_dmac_0_m_dest_axi_araddr
	wire   [2:0] spi_dmac_0_m_dest_axi_arprot;                            // spi_dmac_0:m_dest_axi_arprot -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arprot
	wire  [63:0] spi_dmac_0_m_dest_axi_wdata;                             // spi_dmac_0:m_dest_axi_wdata -> mm_interconnect_1:spi_dmac_0_m_dest_axi_wdata
	wire         spi_dmac_0_m_dest_axi_arvalid;                           // spi_dmac_0:m_dest_axi_arvalid -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arvalid
	wire   [2:0] spi_dmac_0_m_dest_axi_awprot;                            // spi_dmac_0:m_dest_axi_awprot -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awprot
	wire   [3:0] spi_dmac_0_m_dest_axi_awcache;                           // spi_dmac_0:m_dest_axi_awcache -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awcache
	wire         spi_dmac_0_m_dest_axi_arid;                              // spi_dmac_0:m_dest_axi_arid -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arid
	wire   [1:0] spi_dmac_0_m_dest_axi_arlock;                            // spi_dmac_0:m_dest_axi_arlock -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arlock
	wire   [1:0] spi_dmac_0_m_dest_axi_awlock;                            // spi_dmac_0:m_dest_axi_awlock -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awlock
	wire  [31:0] spi_dmac_0_m_dest_axi_awaddr;                            // spi_dmac_0:m_dest_axi_awaddr -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awaddr
	wire   [1:0] spi_dmac_0_m_dest_axi_bresp;                             // mm_interconnect_1:spi_dmac_0_m_dest_axi_bresp -> spi_dmac_0:m_dest_axi_bresp
	wire         spi_dmac_0_m_dest_axi_arready;                           // mm_interconnect_1:spi_dmac_0_m_dest_axi_arready -> spi_dmac_0:m_dest_axi_arready
	wire  [63:0] spi_dmac_0_m_dest_axi_rdata;                             // mm_interconnect_1:spi_dmac_0_m_dest_axi_rdata -> spi_dmac_0:m_dest_axi_rdata
	wire         spi_dmac_0_m_dest_axi_awready;                           // mm_interconnect_1:spi_dmac_0_m_dest_axi_awready -> spi_dmac_0:m_dest_axi_awready
	wire   [1:0] spi_dmac_0_m_dest_axi_arburst;                           // spi_dmac_0:m_dest_axi_arburst -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arburst
	wire   [2:0] spi_dmac_0_m_dest_axi_arsize;                            // spi_dmac_0:m_dest_axi_arsize -> mm_interconnect_1:spi_dmac_0_m_dest_axi_arsize
	wire         spi_dmac_0_m_dest_axi_bready;                            // spi_dmac_0:m_dest_axi_bready -> mm_interconnect_1:spi_dmac_0_m_dest_axi_bready
	wire         spi_dmac_0_m_dest_axi_rlast;                             // mm_interconnect_1:spi_dmac_0_m_dest_axi_rlast -> spi_dmac_0:m_dest_axi_rlast
	wire         spi_dmac_0_m_dest_axi_wlast;                             // spi_dmac_0:m_dest_axi_wlast -> mm_interconnect_1:spi_dmac_0_m_dest_axi_wlast
	wire   [1:0] spi_dmac_0_m_dest_axi_rresp;                             // mm_interconnect_1:spi_dmac_0_m_dest_axi_rresp -> spi_dmac_0:m_dest_axi_rresp
	wire         spi_dmac_0_m_dest_axi_awid;                              // spi_dmac_0:m_dest_axi_awid -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awid
	wire         spi_dmac_0_m_dest_axi_bid;                               // mm_interconnect_1:spi_dmac_0_m_dest_axi_bid -> spi_dmac_0:m_dest_axi_bid
	wire         spi_dmac_0_m_dest_axi_bvalid;                            // mm_interconnect_1:spi_dmac_0_m_dest_axi_bvalid -> spi_dmac_0:m_dest_axi_bvalid
	wire         spi_dmac_0_m_dest_axi_awvalid;                           // spi_dmac_0:m_dest_axi_awvalid -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awvalid
	wire         spi_dmac_0_m_dest_axi_rvalid;                            // mm_interconnect_1:spi_dmac_0_m_dest_axi_rvalid -> spi_dmac_0:m_dest_axi_rvalid
	wire   [2:0] spi_dmac_0_m_dest_axi_awsize;                            // spi_dmac_0:m_dest_axi_awsize -> mm_interconnect_1:spi_dmac_0_m_dest_axi_awsize
	wire   [1:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awburst;       // mm_interconnect_1:sys_hps_f2h_sdram1_data_awburst -> sys_hps:f2h_sdram1_AWBURST
	wire   [3:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_arlen;         // mm_interconnect_1:sys_hps_f2h_sdram1_data_arlen -> sys_hps:f2h_sdram1_ARLEN
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_wstrb;         // mm_interconnect_1:sys_hps_f2h_sdram1_data_wstrb -> sys_hps:f2h_sdram1_WSTRB
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_wready;        // sys_hps:f2h_sdram1_WREADY -> mm_interconnect_1:sys_hps_f2h_sdram1_data_wready
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_rid;           // sys_hps:f2h_sdram1_RID -> mm_interconnect_1:sys_hps_f2h_sdram1_data_rid
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_rready;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_rready -> sys_hps:f2h_sdram1_RREADY
	wire   [3:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awlen;         // mm_interconnect_1:sys_hps_f2h_sdram1_data_awlen -> sys_hps:f2h_sdram1_AWLEN
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_wid;           // mm_interconnect_1:sys_hps_f2h_sdram1_data_wid -> sys_hps:f2h_sdram1_WID
	wire   [3:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_arcache;       // mm_interconnect_1:sys_hps_f2h_sdram1_data_arcache -> sys_hps:f2h_sdram1_ARCACHE
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_wvalid;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_wvalid -> sys_hps:f2h_sdram1_WVALID
	wire  [31:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_araddr;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_araddr -> sys_hps:f2h_sdram1_ARADDR
	wire   [2:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_arprot;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_arprot -> sys_hps:f2h_sdram1_ARPROT
	wire   [2:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awprot;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_awprot -> sys_hps:f2h_sdram1_AWPROT
	wire  [63:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_wdata;         // mm_interconnect_1:sys_hps_f2h_sdram1_data_wdata -> sys_hps:f2h_sdram1_WDATA
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_arvalid;       // mm_interconnect_1:sys_hps_f2h_sdram1_data_arvalid -> sys_hps:f2h_sdram1_ARVALID
	wire   [3:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awcache;       // mm_interconnect_1:sys_hps_f2h_sdram1_data_awcache -> sys_hps:f2h_sdram1_AWCACHE
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_arid;          // mm_interconnect_1:sys_hps_f2h_sdram1_data_arid -> sys_hps:f2h_sdram1_ARID
	wire   [1:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_arlock;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_arlock -> sys_hps:f2h_sdram1_ARLOCK
	wire   [1:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awlock;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_awlock -> sys_hps:f2h_sdram1_AWLOCK
	wire  [31:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awaddr;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_awaddr -> sys_hps:f2h_sdram1_AWADDR
	wire   [1:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_bresp;         // sys_hps:f2h_sdram1_BRESP -> mm_interconnect_1:sys_hps_f2h_sdram1_data_bresp
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_arready;       // sys_hps:f2h_sdram1_ARREADY -> mm_interconnect_1:sys_hps_f2h_sdram1_data_arready
	wire  [63:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_rdata;         // sys_hps:f2h_sdram1_RDATA -> mm_interconnect_1:sys_hps_f2h_sdram1_data_rdata
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_awready;       // sys_hps:f2h_sdram1_AWREADY -> mm_interconnect_1:sys_hps_f2h_sdram1_data_awready
	wire   [1:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_arburst;       // mm_interconnect_1:sys_hps_f2h_sdram1_data_arburst -> sys_hps:f2h_sdram1_ARBURST
	wire   [2:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_arsize;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_arsize -> sys_hps:f2h_sdram1_ARSIZE
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_bready;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_bready -> sys_hps:f2h_sdram1_BREADY
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_rlast;         // sys_hps:f2h_sdram1_RLAST -> mm_interconnect_1:sys_hps_f2h_sdram1_data_rlast
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_wlast;         // mm_interconnect_1:sys_hps_f2h_sdram1_data_wlast -> sys_hps:f2h_sdram1_WLAST
	wire   [1:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_rresp;         // sys_hps:f2h_sdram1_RRESP -> mm_interconnect_1:sys_hps_f2h_sdram1_data_rresp
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awid;          // mm_interconnect_1:sys_hps_f2h_sdram1_data_awid -> sys_hps:f2h_sdram1_AWID
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_bid;           // sys_hps:f2h_sdram1_BID -> mm_interconnect_1:sys_hps_f2h_sdram1_data_bid
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_bvalid;        // sys_hps:f2h_sdram1_BVALID -> mm_interconnect_1:sys_hps_f2h_sdram1_data_bvalid
	wire   [2:0] mm_interconnect_1_sys_hps_f2h_sdram1_data_awsize;        // mm_interconnect_1:sys_hps_f2h_sdram1_data_awsize -> sys_hps:f2h_sdram1_AWSIZE
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_awvalid;       // mm_interconnect_1:sys_hps_f2h_sdram1_data_awvalid -> sys_hps:f2h_sdram1_AWVALID
	wire         mm_interconnect_1_sys_hps_f2h_sdram1_data_rvalid;        // sys_hps:f2h_sdram1_RVALID -> mm_interconnect_1:sys_hps_f2h_sdram1_data_rvalid
	wire   [1:0] hdmi_dmac_0_m_src_axi_awburst;                           // hdmi_dmac_0:m_src_axi_awburst -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awburst
	wire   [3:0] hdmi_dmac_0_m_src_axi_arlen;                             // hdmi_dmac_0:m_src_axi_arlen -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arlen
	wire   [7:0] hdmi_dmac_0_m_src_axi_wstrb;                             // hdmi_dmac_0:m_src_axi_wstrb -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_wstrb
	wire         hdmi_dmac_0_m_src_axi_wready;                            // mm_interconnect_2:hdmi_dmac_0_m_src_axi_wready -> hdmi_dmac_0:m_src_axi_wready
	wire         hdmi_dmac_0_m_src_axi_rid;                               // mm_interconnect_2:hdmi_dmac_0_m_src_axi_rid -> hdmi_dmac_0:m_src_axi_rid
	wire         hdmi_dmac_0_m_src_axi_rready;                            // hdmi_dmac_0:m_src_axi_rready -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_rready
	wire   [3:0] hdmi_dmac_0_m_src_axi_awlen;                             // hdmi_dmac_0:m_src_axi_awlen -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awlen
	wire         hdmi_dmac_0_m_src_axi_wid;                               // hdmi_dmac_0:m_src_axi_wid -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_wid
	wire   [3:0] hdmi_dmac_0_m_src_axi_arcache;                           // hdmi_dmac_0:m_src_axi_arcache -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arcache
	wire         hdmi_dmac_0_m_src_axi_wvalid;                            // hdmi_dmac_0:m_src_axi_wvalid -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_wvalid
	wire  [31:0] hdmi_dmac_0_m_src_axi_araddr;                            // hdmi_dmac_0:m_src_axi_araddr -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_araddr
	wire   [2:0] hdmi_dmac_0_m_src_axi_arprot;                            // hdmi_dmac_0:m_src_axi_arprot -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arprot
	wire  [63:0] hdmi_dmac_0_m_src_axi_wdata;                             // hdmi_dmac_0:m_src_axi_wdata -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_wdata
	wire         hdmi_dmac_0_m_src_axi_arvalid;                           // hdmi_dmac_0:m_src_axi_arvalid -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arvalid
	wire   [2:0] hdmi_dmac_0_m_src_axi_awprot;                            // hdmi_dmac_0:m_src_axi_awprot -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awprot
	wire   [3:0] hdmi_dmac_0_m_src_axi_awcache;                           // hdmi_dmac_0:m_src_axi_awcache -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awcache
	wire         hdmi_dmac_0_m_src_axi_arid;                              // hdmi_dmac_0:m_src_axi_arid -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arid
	wire   [1:0] hdmi_dmac_0_m_src_axi_arlock;                            // hdmi_dmac_0:m_src_axi_arlock -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arlock
	wire   [1:0] hdmi_dmac_0_m_src_axi_awlock;                            // hdmi_dmac_0:m_src_axi_awlock -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awlock
	wire  [31:0] hdmi_dmac_0_m_src_axi_awaddr;                            // hdmi_dmac_0:m_src_axi_awaddr -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awaddr
	wire   [1:0] hdmi_dmac_0_m_src_axi_bresp;                             // mm_interconnect_2:hdmi_dmac_0_m_src_axi_bresp -> hdmi_dmac_0:m_src_axi_bresp
	wire         hdmi_dmac_0_m_src_axi_arready;                           // mm_interconnect_2:hdmi_dmac_0_m_src_axi_arready -> hdmi_dmac_0:m_src_axi_arready
	wire  [63:0] hdmi_dmac_0_m_src_axi_rdata;                             // mm_interconnect_2:hdmi_dmac_0_m_src_axi_rdata -> hdmi_dmac_0:m_src_axi_rdata
	wire         hdmi_dmac_0_m_src_axi_awready;                           // mm_interconnect_2:hdmi_dmac_0_m_src_axi_awready -> hdmi_dmac_0:m_src_axi_awready
	wire   [1:0] hdmi_dmac_0_m_src_axi_arburst;                           // hdmi_dmac_0:m_src_axi_arburst -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arburst
	wire   [2:0] hdmi_dmac_0_m_src_axi_arsize;                            // hdmi_dmac_0:m_src_axi_arsize -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_arsize
	wire         hdmi_dmac_0_m_src_axi_bready;                            // hdmi_dmac_0:m_src_axi_bready -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_bready
	wire         hdmi_dmac_0_m_src_axi_rlast;                             // mm_interconnect_2:hdmi_dmac_0_m_src_axi_rlast -> hdmi_dmac_0:m_src_axi_rlast
	wire         hdmi_dmac_0_m_src_axi_wlast;                             // hdmi_dmac_0:m_src_axi_wlast -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_wlast
	wire   [1:0] hdmi_dmac_0_m_src_axi_rresp;                             // mm_interconnect_2:hdmi_dmac_0_m_src_axi_rresp -> hdmi_dmac_0:m_src_axi_rresp
	wire         hdmi_dmac_0_m_src_axi_awid;                              // hdmi_dmac_0:m_src_axi_awid -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awid
	wire         hdmi_dmac_0_m_src_axi_bid;                               // mm_interconnect_2:hdmi_dmac_0_m_src_axi_bid -> hdmi_dmac_0:m_src_axi_bid
	wire         hdmi_dmac_0_m_src_axi_bvalid;                            // mm_interconnect_2:hdmi_dmac_0_m_src_axi_bvalid -> hdmi_dmac_0:m_src_axi_bvalid
	wire         hdmi_dmac_0_m_src_axi_awvalid;                           // hdmi_dmac_0:m_src_axi_awvalid -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awvalid
	wire         hdmi_dmac_0_m_src_axi_rvalid;                            // mm_interconnect_2:hdmi_dmac_0_m_src_axi_rvalid -> hdmi_dmac_0:m_src_axi_rvalid
	wire   [2:0] hdmi_dmac_0_m_src_axi_awsize;                            // hdmi_dmac_0:m_src_axi_awsize -> mm_interconnect_2:hdmi_dmac_0_m_src_axi_awsize
	wire  [63:0] mm_interconnect_2_sys_hps_f2h_sdram0_data_readdata;      // sys_hps:f2h_sdram0_READDATA -> mm_interconnect_2:sys_hps_f2h_sdram0_data_readdata
	wire         mm_interconnect_2_sys_hps_f2h_sdram0_data_waitrequest;   // sys_hps:f2h_sdram0_WAITREQUEST -> mm_interconnect_2:sys_hps_f2h_sdram0_data_waitrequest
	wire  [28:0] mm_interconnect_2_sys_hps_f2h_sdram0_data_address;       // mm_interconnect_2:sys_hps_f2h_sdram0_data_address -> sys_hps:f2h_sdram0_ADDRESS
	wire         mm_interconnect_2_sys_hps_f2h_sdram0_data_read;          // mm_interconnect_2:sys_hps_f2h_sdram0_data_read -> sys_hps:f2h_sdram0_READ
	wire   [7:0] mm_interconnect_2_sys_hps_f2h_sdram0_data_byteenable;    // mm_interconnect_2:sys_hps_f2h_sdram0_data_byteenable -> sys_hps:f2h_sdram0_BYTEENABLE
	wire         mm_interconnect_2_sys_hps_f2h_sdram0_data_readdatavalid; // sys_hps:f2h_sdram0_READDATAVALID -> mm_interconnect_2:sys_hps_f2h_sdram0_data_readdatavalid
	wire         mm_interconnect_2_sys_hps_f2h_sdram0_data_write;         // mm_interconnect_2:sys_hps_f2h_sdram0_data_write -> sys_hps:f2h_sdram0_WRITE
	wire  [63:0] mm_interconnect_2_sys_hps_f2h_sdram0_data_writedata;     // mm_interconnect_2:sys_hps_f2h_sdram0_data_writedata -> sys_hps:f2h_sdram0_WRITEDATA
	wire   [7:0] mm_interconnect_2_sys_hps_f2h_sdram0_data_burstcount;    // mm_interconnect_2:sys_hps_f2h_sdram0_data_burstcount -> sys_hps:f2h_sdram0_BURSTCOUNT
	wire         irq_mapper_receiver0_irq;                                // hdmi_dmac_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                // spi_dmac_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                // sys_gpio_bd:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                // sys_gpio_in:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                // axi_spi_engine_0:irq -> irq_mapper:receiver4_irq
	wire  [31:0] sys_hps_f2h_irq0_irq;                                    // irq_mapper:sender_irq -> sys_hps:f2h_irq_p0
	wire  [31:0] sys_hps_f2h_irq1_irq;                                    // irq_mapper_001:sender_irq -> sys_hps:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [axi_hdmi_tx_0:s_axi_aresetn, axi_spi_engine_0:s_axi_aresetn, hdmi_dmac_0:m_src_axi_aresetn, hdmi_dmac_0:s_axi_aresetn, mm_interconnect_0:sys_id_reset_reset_bridge_in_reset_reset, mm_interconnect_1:spi_dmac_0_m_dest_axi_reset_reset_bridge_in_reset_reset, mm_interconnect_2:hdmi_dmac_0_m_src_axi_reset_reset_bridge_in_reset_reset, spi_dmac_0:m_dest_axi_aresetn, spi_dmac_0:s_axi_aresetn, sys_gpio_bd:reset_n, sys_gpio_in:reset_n, sys_gpio_out:reset_n, sys_id:reset_n]
	wire         rst_controller_001_reset_out_reset;                      // rst_controller_001:reset_out -> [mm_interconnect_0:sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:spi_dmac_0_m_dest_axi_id_pad_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sys_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset]

	axi_hdmi_tx #(
		.ID               (0),
		.FPGA_TECHNOLOGY  (101),
		.INTERFACE        ("16_BIT"),
		.CR_CB_N          (0),
		.OUT_CLK_POLARITY (0)
	) axi_hdmi_tx_0 (
		.s_axi_aclk        (sys_hps_h2f_user1_clock_clk),                   // s_axi_clock.clk
		.s_axi_awvalid     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awvalid), //       s_axi.awvalid
		.s_axi_awaddr      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awaddr),  //            .awaddr
		.s_axi_awprot      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awprot),  //            .awprot
		.s_axi_awready     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awready), //            .awready
		.s_axi_wvalid      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wvalid),  //            .wvalid
		.s_axi_wdata       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wdata),   //            .wdata
		.s_axi_wstrb       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wstrb),   //            .wstrb
		.s_axi_wready      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wready),  //            .wready
		.s_axi_bvalid      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bvalid),  //            .bvalid
		.s_axi_bresp       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bresp),   //            .bresp
		.s_axi_bready      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bready),  //            .bready
		.s_axi_arvalid     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arvalid), //            .arvalid
		.s_axi_araddr      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_araddr),  //            .araddr
		.s_axi_arprot      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arprot),  //            .arprot
		.s_axi_arready     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arready), //            .arready
		.s_axi_rvalid      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rvalid),  //            .rvalid
		.s_axi_rresp       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rresp),   //            .rresp
		.s_axi_rdata       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rdata),   //            .rdata
		.s_axi_rready      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rready),  //            .rready
		.hdmi_clk          (hdmi_pll_outclk0_clk),                          //  hdmi_clock.clk
		.hdmi_out_clk      (hdmi_out_h_clk),                                //     hdmi_if.h_clk
		.hdmi_16_hsync     (hdmi_out_h16_hsync),                            //            .h16_hsync
		.hdmi_16_vsync     (hdmi_out_h16_vsync),                            //            .h16_vsync
		.hdmi_16_data_e    (hdmi_out_h16_data_e),                           //            .h16_data_e
		.hdmi_16_data      (hdmi_out_h16_data),                             //            .h16_data
		.hdmi_16_es_data   (hdmi_out_h16_es_data),                          //            .h16_es_data
		.hdmi_24_hsync     (hdmi_out_h24_hsync),                            //            .h24_hsync
		.hdmi_24_vsync     (hdmi_out_h24_vsync),                            //            .h24_vsync
		.hdmi_24_data_e    (hdmi_out_h24_data_e),                           //            .h24_data_e
		.hdmi_24_data      (hdmi_out_h24_data),                             //            .h24_data
		.hdmi_36_hsync     (hdmi_out_h36_hsync),                            //            .h36_hsync
		.hdmi_36_vsync     (hdmi_out_h36_vsync),                            //            .h36_vsync
		.hdmi_36_data_e    (hdmi_out_h36_data_e),                           //            .h36_data_e
		.hdmi_36_data      (hdmi_out_h36_data),                             //            .h36_data
		.vdma_clk          (sys_hps_h2f_user1_clock_clk),                   //  vdma_clock.clk
		.s_axi_aresetn     (~rst_controller_reset_out_reset),               //  vdma_reset.reset_n
		.vdma_end_of_frame (hdmi_dmac_0_m_axis_tlast),                      //     vdma_if.tlast
		.vdma_valid        (hdmi_dmac_0_m_axis_tvalid),                     //            .tvalid
		.vdma_data         (hdmi_dmac_0_m_axis_tdata),                      //            .tdata
		.vdma_ready        (hdmi_dmac_0_m_axis_tready)                      //            .tready
	);

	axi_spi_engine #(
		.CMD_FIFO_ADDRESS_WIDTH         (4),
		.SYNC_FIFO_ADDRESS_WIDTH        (4),
		.SDO_FIFO_ADDRESS_WIDTH         (5),
		.SDI_FIFO_ADDRESS_WIDTH         (5),
		.MM_IF_TYPE                     (0),
		.ASYNC_SPI_CLK                  (1),
		.NUM_OFFLOAD                    (1),
		.OFFLOAD0_CMD_MEM_ADDRESS_WIDTH (4),
		.OFFLOAD0_SDO_MEM_ADDRESS_WIDTH (4),
		.ID                             (0),
		.DATA_WIDTH                     (18),
		.NUM_OF_SDI                     (2)
	) axi_spi_engine_0 (
		.s_axi_aclk           (sys_hps_h2f_user1_clock_clk),                           //               s_axi_aclk.clk
		.s_axi_aresetn        (~rst_controller_reset_out_reset),                       //            s_axi_aresetn.reset_n
		.s_axi_awvalid        (mm_interconnect_0_axi_spi_engine_0_s_axi_awvalid),      //                    s_axi.awvalid
		.s_axi_awaddr         (mm_interconnect_0_axi_spi_engine_0_s_axi_awaddr),       //                         .awaddr
		.s_axi_awready        (mm_interconnect_0_axi_spi_engine_0_s_axi_awready),      //                         .awready
		.s_axi_awprot         (mm_interconnect_0_axi_spi_engine_0_s_axi_awprot),       //                         .awprot
		.s_axi_wvalid         (mm_interconnect_0_axi_spi_engine_0_s_axi_wvalid),       //                         .wvalid
		.s_axi_wdata          (mm_interconnect_0_axi_spi_engine_0_s_axi_wdata),        //                         .wdata
		.s_axi_wstrb          (mm_interconnect_0_axi_spi_engine_0_s_axi_wstrb),        //                         .wstrb
		.s_axi_wready         (mm_interconnect_0_axi_spi_engine_0_s_axi_wready),       //                         .wready
		.s_axi_bvalid         (mm_interconnect_0_axi_spi_engine_0_s_axi_bvalid),       //                         .bvalid
		.s_axi_bresp          (mm_interconnect_0_axi_spi_engine_0_s_axi_bresp),        //                         .bresp
		.s_axi_bready         (mm_interconnect_0_axi_spi_engine_0_s_axi_bready),       //                         .bready
		.s_axi_arvalid        (mm_interconnect_0_axi_spi_engine_0_s_axi_arvalid),      //                         .arvalid
		.s_axi_araddr         (mm_interconnect_0_axi_spi_engine_0_s_axi_araddr),       //                         .araddr
		.s_axi_arready        (mm_interconnect_0_axi_spi_engine_0_s_axi_arready),      //                         .arready
		.s_axi_arprot         (mm_interconnect_0_axi_spi_engine_0_s_axi_arprot),       //                         .arprot
		.s_axi_rvalid         (mm_interconnect_0_axi_spi_engine_0_s_axi_rvalid),       //                         .rvalid
		.s_axi_rready         (mm_interconnect_0_axi_spi_engine_0_s_axi_rready),       //                         .rready
		.s_axi_rresp          (mm_interconnect_0_axi_spi_engine_0_s_axi_rresp),        //                         .rresp
		.s_axi_rdata          (mm_interconnect_0_axi_spi_engine_0_s_axi_rdata),        //                         .rdata
		.spi_clk              (spi_engine_pll_outclk0_clk),                            //                  spi_clk.clk
		.spi_resetn           (axi_spi_engine_0_spi_resetn_reset),                     //               spi_resetn.reset_n
		.cmd_ready            (spi_engine_interconnect_0_s1_ctrl_cmd_ready),           //          spi_engine_ctrl.cmd_ready
		.cmd_valid            (axi_spi_engine_0_spi_engine_ctrl_cmd_valid),            //                         .cmd_valid
		.cmd_data             (axi_spi_engine_0_spi_engine_ctrl_cmd_data),             //                         .cmd_data
		.sdo_data_ready       (spi_engine_interconnect_0_s1_ctrl_sdo_ready),           //                         .sdo_ready
		.sdo_data_valid       (axi_spi_engine_0_spi_engine_ctrl_sdo_valid),            //                         .sdo_valid
		.sdo_data             (axi_spi_engine_0_spi_engine_ctrl_sdo_data),             //                         .sdo_data
		.sdi_data_ready       (axi_spi_engine_0_spi_engine_ctrl_sdi_ready),            //                         .sdi_ready
		.sdi_data_valid       (spi_engine_interconnect_0_s1_ctrl_sdi_valid),           //                         .sdi_valid
		.sdi_data             (spi_engine_interconnect_0_s1_ctrl_sdi_data),            //                         .sdi_data
		.sync_ready           (axi_spi_engine_0_spi_engine_ctrl_sync_ready),           //                         .sync_ready
		.sync_valid           (spi_engine_interconnect_0_s1_ctrl_sync_valid),          //                         .sync_valid
		.sync_data            (spi_engine_interconnect_0_s1_ctrl_sync_data),           //                         .sync_data
		.offload0_cmd_wr_en   (axi_spi_engine_0_spi_engine_offload_ctrl0_cmd_wr_en),   // spi_engine_offload_ctrl0.cmd_wr_en
		.offload0_cmd_wr_data (axi_spi_engine_0_spi_engine_offload_ctrl0_cmd_wr_data), //                         .cmd_wr_data
		.offload0_sdo_wr_en   (axi_spi_engine_0_spi_engine_offload_ctrl0_sdo_wr_en),   //                         .sdo_wr_en
		.offload0_sdo_wr_data (axi_spi_engine_0_spi_engine_offload_ctrl0_sdo_wr_data), //                         .sdo_wr_data
		.offload0_mem_reset   (axi_spi_engine_0_spi_engine_offload_ctrl0_reset),       //                         .reset
		.offload0_enable      (axi_spi_engine_0_spi_engine_offload_ctrl0_enable),      //                         .enable
		.offload0_enabled     (spi_engine_offload_0_spi_engine_offload_ctrl_enabled),  //                         .enabled
		.irq                  (irq_mapper_receiver4_irq),                              //                      irq.irq
		.pulse_gen_period     (),                                                      //         pulse_gen_period.pulse_gen_period
		.pulse_gen_load       ()                                                       //           pulse_gen_load.pulse_gen_load
	);

	axi_dmac #(
		.ID                    (0),
		.DMA_LENGTH_WIDTH      (24),
		.FIFO_SIZE             (8),
		.MAX_BYTES_PER_BURST   (128),
		.DMA_TYPE_SRC          (0),
		.DMA_AXI_PROTOCOL_SRC  (1),
		.DMA_DATA_WIDTH_SRC    (64),
		.AXI_SLICE_SRC         (0),
		.DMA_TYPE_DEST         (1),
		.DMA_AXI_PROTOCOL_DEST (1),
		.DMA_DATA_WIDTH_DEST   (64),
		.AXI_SLICE_DEST        (0),
		.CYCLIC                (1),
		.DMA_2D_TRANSFER       (1),
		.SYNC_TRANSFER_START   (0),
		.ASYNC_CLK_REQ_SRC     (0),
		.ASYNC_CLK_SRC_DEST    (0),
		.ASYNC_CLK_DEST_REQ    (0),
		.ENABLE_DIAGNOSTICS_IF (0),
		.DMA_AXIS_ID_W         (8),
		.DMA_AXIS_DEST_W       (4)
	) hdmi_dmac_0 (
		.s_axi_aclk             (sys_hps_h2f_user1_clock_clk),                                          //        s_axi_clock.clk
		.s_axi_aresetn          (~rst_controller_reset_out_reset),                                      //        s_axi_reset.reset_n
		.s_axi_awvalid          (mm_interconnect_0_hdmi_dmac_0_s_axi_awvalid),                          //              s_axi.awvalid
		.s_axi_awaddr           (mm_interconnect_0_hdmi_dmac_0_s_axi_awaddr),                           //                   .awaddr
		.s_axi_awprot           (mm_interconnect_0_hdmi_dmac_0_s_axi_awprot),                           //                   .awprot
		.s_axi_awready          (mm_interconnect_0_hdmi_dmac_0_s_axi_awready),                          //                   .awready
		.s_axi_wvalid           (mm_interconnect_0_hdmi_dmac_0_s_axi_wvalid),                           //                   .wvalid
		.s_axi_wdata            (mm_interconnect_0_hdmi_dmac_0_s_axi_wdata),                            //                   .wdata
		.s_axi_wstrb            (mm_interconnect_0_hdmi_dmac_0_s_axi_wstrb),                            //                   .wstrb
		.s_axi_wready           (mm_interconnect_0_hdmi_dmac_0_s_axi_wready),                           //                   .wready
		.s_axi_bvalid           (mm_interconnect_0_hdmi_dmac_0_s_axi_bvalid),                           //                   .bvalid
		.s_axi_bresp            (mm_interconnect_0_hdmi_dmac_0_s_axi_bresp),                            //                   .bresp
		.s_axi_bready           (mm_interconnect_0_hdmi_dmac_0_s_axi_bready),                           //                   .bready
		.s_axi_arvalid          (mm_interconnect_0_hdmi_dmac_0_s_axi_arvalid),                          //                   .arvalid
		.s_axi_araddr           (mm_interconnect_0_hdmi_dmac_0_s_axi_araddr),                           //                   .araddr
		.s_axi_arprot           (mm_interconnect_0_hdmi_dmac_0_s_axi_arprot),                           //                   .arprot
		.s_axi_arready          (mm_interconnect_0_hdmi_dmac_0_s_axi_arready),                          //                   .arready
		.s_axi_rvalid           (mm_interconnect_0_hdmi_dmac_0_s_axi_rvalid),                           //                   .rvalid
		.s_axi_rresp            (mm_interconnect_0_hdmi_dmac_0_s_axi_rresp),                            //                   .rresp
		.s_axi_rdata            (mm_interconnect_0_hdmi_dmac_0_s_axi_rdata),                            //                   .rdata
		.s_axi_rready           (mm_interconnect_0_hdmi_dmac_0_s_axi_rready),                           //                   .rready
		.irq                    (irq_mapper_receiver0_irq),                                             //   interrupt_sender.irq
		.m_src_axi_aclk         (sys_hps_h2f_user1_clock_clk),                                          //    m_src_axi_clock.clk
		.m_src_axi_aresetn      (~rst_controller_reset_out_reset),                                      //    m_src_axi_reset.reset_n
		.m_axis_aclk            (sys_hps_h2f_user1_clock_clk),                                          //     if_m_axis_aclk.clk
		.m_axis_xfer_req        (),                                                                     // if_m_axis_xfer_req.xfer_req
		.m_axis_valid           (hdmi_dmac_0_m_axis_tvalid),                                            //             m_axis.tvalid
		.m_axis_last            (hdmi_dmac_0_m_axis_tlast),                                             //                   .tlast
		.m_axis_ready           (hdmi_dmac_0_m_axis_tready),                                            //                   .tready
		.m_axis_data            (hdmi_dmac_0_m_axis_tdata),                                             //                   .tdata
		.m_src_axi_awvalid      (hdmi_dmac_0_m_src_axi_awvalid),                                        //          m_src_axi.awvalid
		.m_src_axi_awaddr       (hdmi_dmac_0_m_src_axi_awaddr),                                         //                   .awaddr
		.m_src_axi_awready      (hdmi_dmac_0_m_src_axi_awready),                                        //                   .awready
		.m_src_axi_wvalid       (hdmi_dmac_0_m_src_axi_wvalid),                                         //                   .wvalid
		.m_src_axi_wdata        (hdmi_dmac_0_m_src_axi_wdata),                                          //                   .wdata
		.m_src_axi_wstrb        (hdmi_dmac_0_m_src_axi_wstrb),                                          //                   .wstrb
		.m_src_axi_wready       (hdmi_dmac_0_m_src_axi_wready),                                         //                   .wready
		.m_src_axi_bvalid       (hdmi_dmac_0_m_src_axi_bvalid),                                         //                   .bvalid
		.m_src_axi_bresp        (hdmi_dmac_0_m_src_axi_bresp),                                          //                   .bresp
		.m_src_axi_bready       (hdmi_dmac_0_m_src_axi_bready),                                         //                   .bready
		.m_src_axi_arvalid      (hdmi_dmac_0_m_src_axi_arvalid),                                        //                   .arvalid
		.m_src_axi_araddr       (hdmi_dmac_0_m_src_axi_araddr),                                         //                   .araddr
		.m_src_axi_arready      (hdmi_dmac_0_m_src_axi_arready),                                        //                   .arready
		.m_src_axi_rvalid       (hdmi_dmac_0_m_src_axi_rvalid),                                         //                   .rvalid
		.m_src_axi_rresp        (hdmi_dmac_0_m_src_axi_rresp),                                          //                   .rresp
		.m_src_axi_rdata        (hdmi_dmac_0_m_src_axi_rdata),                                          //                   .rdata
		.m_src_axi_rready       (hdmi_dmac_0_m_src_axi_rready),                                         //                   .rready
		.m_src_axi_awlen        (hdmi_dmac_0_m_src_axi_awlen),                                          //                   .awlen
		.m_src_axi_awsize       (hdmi_dmac_0_m_src_axi_awsize),                                         //                   .awsize
		.m_src_axi_awburst      (hdmi_dmac_0_m_src_axi_awburst),                                        //                   .awburst
		.m_src_axi_awcache      (hdmi_dmac_0_m_src_axi_awcache),                                        //                   .awcache
		.m_src_axi_awprot       (hdmi_dmac_0_m_src_axi_awprot),                                         //                   .awprot
		.m_src_axi_wlast        (hdmi_dmac_0_m_src_axi_wlast),                                          //                   .wlast
		.m_src_axi_arlen        (hdmi_dmac_0_m_src_axi_arlen),                                          //                   .arlen
		.m_src_axi_arsize       (hdmi_dmac_0_m_src_axi_arsize),                                         //                   .arsize
		.m_src_axi_arburst      (hdmi_dmac_0_m_src_axi_arburst),                                        //                   .arburst
		.m_src_axi_arcache      (hdmi_dmac_0_m_src_axi_arcache),                                        //                   .arcache
		.m_src_axi_arprot       (hdmi_dmac_0_m_src_axi_arprot),                                         //                   .arprot
		.m_src_axi_awid         (hdmi_dmac_0_m_src_axi_awid),                                           //                   .awid
		.m_src_axi_awlock       (hdmi_dmac_0_m_src_axi_awlock),                                         //                   .awlock
		.m_src_axi_wid          (hdmi_dmac_0_m_src_axi_wid),                                            //                   .wid
		.m_src_axi_arid         (hdmi_dmac_0_m_src_axi_arid),                                           //                   .arid
		.m_src_axi_arlock       (hdmi_dmac_0_m_src_axi_arlock),                                         //                   .arlock
		.m_src_axi_rid          (hdmi_dmac_0_m_src_axi_rid),                                            //                   .rid
		.m_src_axi_bid          (hdmi_dmac_0_m_src_axi_bid),                                            //                   .bid
		.m_src_axi_rlast        (hdmi_dmac_0_m_src_axi_rlast),                                          //                   .rlast
		.m_axis_user            (),                                                                     //        (terminated)
		.m_axis_id              (),                                                                     //        (terminated)
		.m_axis_dest            (),                                                                     //        (terminated)
		.m_axis_strb            (),                                                                     //        (terminated)
		.m_axis_keep            (),                                                                     //        (terminated)
		.m_dest_axi_aclk        (1'b0),                                                                 //        (terminated)
		.m_dest_axi_aresetn     (1'b1),                                                                 //        (terminated)
		.s_axis_aclk            (1'b0),                                                                 //        (terminated)
		.s_axis_xfer_req        (),                                                                     //        (terminated)
		.s_axis_valid           (1'b0),                                                                 //        (terminated)
		.s_axis_last            (1'b0),                                                                 //        (terminated)
		.s_axis_ready           (),                                                                     //        (terminated)
		.s_axis_data            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.s_axis_user            (1'b0),                                                                 //        (terminated)
		.s_axis_id              (8'b00000000),                                                          //        (terminated)
		.s_axis_dest            (4'b0000),                                                              //        (terminated)
		.s_axis_strb            (8'b00000000),                                                          //        (terminated)
		.s_axis_keep            (8'b00000000),                                                          //        (terminated)
		.fifo_rd_clk            (1'b0),                                                                 //        (terminated)
		.fifo_rd_en             (1'b0),                                                                 //        (terminated)
		.fifo_rd_valid          (),                                                                     //        (terminated)
		.fifo_rd_dout           (),                                                                     //        (terminated)
		.fifo_rd_underflow      (),                                                                     //        (terminated)
		.fifo_rd_xfer_req       (),                                                                     //        (terminated)
		.fifo_wr_clk            (1'b0),                                                                 //        (terminated)
		.fifo_wr_en             (1'b0),                                                                 //        (terminated)
		.fifo_wr_din            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.fifo_wr_overflow       (),                                                                     //        (terminated)
		.fifo_wr_sync           (1'b0),                                                                 //        (terminated)
		.fifo_wr_xfer_req       (),                                                                     //        (terminated)
		.dest_diag_level_bursts (),                                                                     //        (terminated)
		.m_dest_axi_awvalid     (),                                                                     //        (terminated)
		.m_dest_axi_awaddr      (),                                                                     //        (terminated)
		.m_dest_axi_awready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_wvalid      (),                                                                     //        (terminated)
		.m_dest_axi_wdata       (),                                                                     //        (terminated)
		.m_dest_axi_wstrb       (),                                                                     //        (terminated)
		.m_dest_axi_wready      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_bready      (),                                                                     //        (terminated)
		.m_dest_axi_arvalid     (),                                                                     //        (terminated)
		.m_dest_axi_araddr      (),                                                                     //        (terminated)
		.m_dest_axi_arready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_rdata       (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.m_dest_axi_rready      (),                                                                     //        (terminated)
		.m_dest_axi_awlen       (),                                                                     //        (terminated)
		.m_dest_axi_awsize      (),                                                                     //        (terminated)
		.m_dest_axi_awburst     (),                                                                     //        (terminated)
		.m_dest_axi_awcache     (),                                                                     //        (terminated)
		.m_dest_axi_awprot      (),                                                                     //        (terminated)
		.m_dest_axi_wlast       (),                                                                     //        (terminated)
		.m_dest_axi_arlen       (),                                                                     //        (terminated)
		.m_dest_axi_arsize      (),                                                                     //        (terminated)
		.m_dest_axi_arburst     (),                                                                     //        (terminated)
		.m_dest_axi_arcache     (),                                                                     //        (terminated)
		.m_dest_axi_arprot      (),                                                                     //        (terminated)
		.m_dest_axi_awid        (),                                                                     //        (terminated)
		.m_dest_axi_awlock      (),                                                                     //        (terminated)
		.m_dest_axi_wid         (),                                                                     //        (terminated)
		.m_dest_axi_arid        (),                                                                     //        (terminated)
		.m_dest_axi_arlock      (),                                                                     //        (terminated)
		.m_dest_axi_rid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rlast       (1'b0)                                                                  //        (terminated)
	);

	system_bd_hdmi_pll hdmi_pll (
		.refclk   (sys_hps_h2f_user1_clock_clk), //  refclk.clk
		.rst      (~sys_rst_reset_n),            //   reset.reset
		.outclk_0 (hdmi_pll_outclk0_clk),        // outclk0.clk
		.locked   ()                             // (terminated)
	);

	axi_dmac #(
		.ID                    (0),
		.DMA_LENGTH_WIDTH      (24),
		.FIFO_SIZE             (8),
		.MAX_BYTES_PER_BURST   (128),
		.DMA_TYPE_SRC          (1),
		.DMA_AXI_PROTOCOL_SRC  (1),
		.DMA_DATA_WIDTH_SRC    (64),
		.AXI_SLICE_SRC         (0),
		.DMA_TYPE_DEST         (0),
		.DMA_AXI_PROTOCOL_DEST (1),
		.DMA_DATA_WIDTH_DEST   (64),
		.AXI_SLICE_DEST        (1),
		.CYCLIC                (0),
		.DMA_2D_TRANSFER       (0),
		.SYNC_TRANSFER_START   (0),
		.ASYNC_CLK_REQ_SRC     (1),
		.ASYNC_CLK_SRC_DEST    (1),
		.ASYNC_CLK_DEST_REQ    (0),
		.ENABLE_DIAGNOSTICS_IF (0),
		.DMA_AXIS_ID_W         (8),
		.DMA_AXIS_DEST_W       (4)
	) spi_dmac_0 (
		.s_axi_aclk             (sys_hps_h2f_user1_clock_clk),                                          //        s_axi_clock.clk
		.s_axi_aresetn          (~rst_controller_reset_out_reset),                                      //        s_axi_reset.reset_n
		.s_axi_awvalid          (mm_interconnect_0_spi_dmac_0_s_axi_awvalid),                           //              s_axi.awvalid
		.s_axi_awaddr           (mm_interconnect_0_spi_dmac_0_s_axi_awaddr),                            //                   .awaddr
		.s_axi_awprot           (mm_interconnect_0_spi_dmac_0_s_axi_awprot),                            //                   .awprot
		.s_axi_awready          (mm_interconnect_0_spi_dmac_0_s_axi_awready),                           //                   .awready
		.s_axi_wvalid           (mm_interconnect_0_spi_dmac_0_s_axi_wvalid),                            //                   .wvalid
		.s_axi_wdata            (mm_interconnect_0_spi_dmac_0_s_axi_wdata),                             //                   .wdata
		.s_axi_wstrb            (mm_interconnect_0_spi_dmac_0_s_axi_wstrb),                             //                   .wstrb
		.s_axi_wready           (mm_interconnect_0_spi_dmac_0_s_axi_wready),                            //                   .wready
		.s_axi_bvalid           (mm_interconnect_0_spi_dmac_0_s_axi_bvalid),                            //                   .bvalid
		.s_axi_bresp            (mm_interconnect_0_spi_dmac_0_s_axi_bresp),                             //                   .bresp
		.s_axi_bready           (mm_interconnect_0_spi_dmac_0_s_axi_bready),                            //                   .bready
		.s_axi_arvalid          (mm_interconnect_0_spi_dmac_0_s_axi_arvalid),                           //                   .arvalid
		.s_axi_araddr           (mm_interconnect_0_spi_dmac_0_s_axi_araddr),                            //                   .araddr
		.s_axi_arprot           (mm_interconnect_0_spi_dmac_0_s_axi_arprot),                            //                   .arprot
		.s_axi_arready          (mm_interconnect_0_spi_dmac_0_s_axi_arready),                           //                   .arready
		.s_axi_rvalid           (mm_interconnect_0_spi_dmac_0_s_axi_rvalid),                            //                   .rvalid
		.s_axi_rresp            (mm_interconnect_0_spi_dmac_0_s_axi_rresp),                             //                   .rresp
		.s_axi_rdata            (mm_interconnect_0_spi_dmac_0_s_axi_rdata),                             //                   .rdata
		.s_axi_rready           (mm_interconnect_0_spi_dmac_0_s_axi_rready),                            //                   .rready
		.irq                    (irq_mapper_receiver1_irq),                                             //   interrupt_sender.irq
		.m_dest_axi_aclk        (sys_hps_h2f_user1_clock_clk),                                          //   m_dest_axi_clock.clk
		.m_dest_axi_aresetn     (~rst_controller_reset_out_reset),                                      //   m_dest_axi_reset.reset_n
		.s_axis_aclk            (spi_engine_pll_outclk0_clk),                                           //     if_s_axis_aclk.clk
		.s_axis_xfer_req        (),                                                                     // if_s_axis_xfer_req.xfer_req
		.s_axis_valid           (upscale_converter_0_m_axis_tvalid),                                    //             s_axis.tvalid
		.s_axis_ready           (upscale_converter_0_m_axis_tready),                                    //                   .tready
		.s_axis_data            (upscale_converter_0_m_axis_tdata),                                     //                   .tdata
		.m_dest_axi_awvalid     (spi_dmac_0_m_dest_axi_awvalid),                                        //         m_dest_axi.awvalid
		.m_dest_axi_awaddr      (spi_dmac_0_m_dest_axi_awaddr),                                         //                   .awaddr
		.m_dest_axi_awready     (spi_dmac_0_m_dest_axi_awready),                                        //                   .awready
		.m_dest_axi_wvalid      (spi_dmac_0_m_dest_axi_wvalid),                                         //                   .wvalid
		.m_dest_axi_wdata       (spi_dmac_0_m_dest_axi_wdata),                                          //                   .wdata
		.m_dest_axi_wstrb       (spi_dmac_0_m_dest_axi_wstrb),                                          //                   .wstrb
		.m_dest_axi_wready      (spi_dmac_0_m_dest_axi_wready),                                         //                   .wready
		.m_dest_axi_bvalid      (spi_dmac_0_m_dest_axi_bvalid),                                         //                   .bvalid
		.m_dest_axi_bresp       (spi_dmac_0_m_dest_axi_bresp),                                          //                   .bresp
		.m_dest_axi_bready      (spi_dmac_0_m_dest_axi_bready),                                         //                   .bready
		.m_dest_axi_arvalid     (spi_dmac_0_m_dest_axi_arvalid),                                        //                   .arvalid
		.m_dest_axi_araddr      (spi_dmac_0_m_dest_axi_araddr),                                         //                   .araddr
		.m_dest_axi_arready     (spi_dmac_0_m_dest_axi_arready),                                        //                   .arready
		.m_dest_axi_rvalid      (spi_dmac_0_m_dest_axi_rvalid),                                         //                   .rvalid
		.m_dest_axi_rresp       (spi_dmac_0_m_dest_axi_rresp),                                          //                   .rresp
		.m_dest_axi_rdata       (spi_dmac_0_m_dest_axi_rdata),                                          //                   .rdata
		.m_dest_axi_rready      (spi_dmac_0_m_dest_axi_rready),                                         //                   .rready
		.m_dest_axi_awlen       (spi_dmac_0_m_dest_axi_awlen),                                          //                   .awlen
		.m_dest_axi_awsize      (spi_dmac_0_m_dest_axi_awsize),                                         //                   .awsize
		.m_dest_axi_awburst     (spi_dmac_0_m_dest_axi_awburst),                                        //                   .awburst
		.m_dest_axi_awcache     (spi_dmac_0_m_dest_axi_awcache),                                        //                   .awcache
		.m_dest_axi_awprot      (spi_dmac_0_m_dest_axi_awprot),                                         //                   .awprot
		.m_dest_axi_wlast       (spi_dmac_0_m_dest_axi_wlast),                                          //                   .wlast
		.m_dest_axi_arlen       (spi_dmac_0_m_dest_axi_arlen),                                          //                   .arlen
		.m_dest_axi_arsize      (spi_dmac_0_m_dest_axi_arsize),                                         //                   .arsize
		.m_dest_axi_arburst     (spi_dmac_0_m_dest_axi_arburst),                                        //                   .arburst
		.m_dest_axi_arcache     (spi_dmac_0_m_dest_axi_arcache),                                        //                   .arcache
		.m_dest_axi_arprot      (spi_dmac_0_m_dest_axi_arprot),                                         //                   .arprot
		.m_dest_axi_awid        (spi_dmac_0_m_dest_axi_awid),                                           //                   .awid
		.m_dest_axi_awlock      (spi_dmac_0_m_dest_axi_awlock),                                         //                   .awlock
		.m_dest_axi_wid         (spi_dmac_0_m_dest_axi_wid),                                            //                   .wid
		.m_dest_axi_arid        (spi_dmac_0_m_dest_axi_arid),                                           //                   .arid
		.m_dest_axi_arlock      (spi_dmac_0_m_dest_axi_arlock),                                         //                   .arlock
		.m_dest_axi_rid         (spi_dmac_0_m_dest_axi_rid),                                            //                   .rid
		.m_dest_axi_bid         (spi_dmac_0_m_dest_axi_bid),                                            //                   .bid
		.m_dest_axi_rlast       (spi_dmac_0_m_dest_axi_rlast),                                          //                   .rlast
		.s_axis_last            (1'b0),                                                                 //        (terminated)
		.s_axis_user            (1'b0),                                                                 //        (terminated)
		.s_axis_id              (8'b00000000),                                                          //        (terminated)
		.s_axis_dest            (4'b0000),                                                              //        (terminated)
		.s_axis_strb            (8'b11111111),                                                          //        (terminated)
		.s_axis_keep            (8'b11111111),                                                          //        (terminated)
		.m_src_axi_aclk         (1'b0),                                                                 //        (terminated)
		.m_src_axi_aresetn      (1'b1),                                                                 //        (terminated)
		.m_axis_aclk            (1'b0),                                                                 //        (terminated)
		.m_axis_xfer_req        (),                                                                     //        (terminated)
		.m_axis_valid           (),                                                                     //        (terminated)
		.m_axis_last            (),                                                                     //        (terminated)
		.m_axis_ready           (1'b0),                                                                 //        (terminated)
		.m_axis_data            (),                                                                     //        (terminated)
		.m_axis_user            (),                                                                     //        (terminated)
		.m_axis_id              (),                                                                     //        (terminated)
		.m_axis_dest            (),                                                                     //        (terminated)
		.m_axis_strb            (),                                                                     //        (terminated)
		.m_axis_keep            (),                                                                     //        (terminated)
		.fifo_rd_clk            (1'b0),                                                                 //        (terminated)
		.fifo_rd_en             (1'b0),                                                                 //        (terminated)
		.fifo_rd_valid          (),                                                                     //        (terminated)
		.fifo_rd_dout           (),                                                                     //        (terminated)
		.fifo_rd_underflow      (),                                                                     //        (terminated)
		.fifo_rd_xfer_req       (),                                                                     //        (terminated)
		.fifo_wr_clk            (1'b0),                                                                 //        (terminated)
		.fifo_wr_en             (1'b0),                                                                 //        (terminated)
		.fifo_wr_din            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.fifo_wr_overflow       (),                                                                     //        (terminated)
		.fifo_wr_sync           (1'b0),                                                                 //        (terminated)
		.fifo_wr_xfer_req       (),                                                                     //        (terminated)
		.dest_diag_level_bursts (),                                                                     //        (terminated)
		.m_src_axi_awvalid      (),                                                                     //        (terminated)
		.m_src_axi_awaddr       (),                                                                     //        (terminated)
		.m_src_axi_awready      (1'b0),                                                                 //        (terminated)
		.m_src_axi_wvalid       (),                                                                     //        (terminated)
		.m_src_axi_wdata        (),                                                                     //        (terminated)
		.m_src_axi_wstrb        (),                                                                     //        (terminated)
		.m_src_axi_wready       (1'b0),                                                                 //        (terminated)
		.m_src_axi_bvalid       (1'b0),                                                                 //        (terminated)
		.m_src_axi_bresp        (2'b00),                                                                //        (terminated)
		.m_src_axi_bready       (),                                                                     //        (terminated)
		.m_src_axi_arvalid      (),                                                                     //        (terminated)
		.m_src_axi_araddr       (),                                                                     //        (terminated)
		.m_src_axi_arready      (1'b0),                                                                 //        (terminated)
		.m_src_axi_rvalid       (1'b0),                                                                 //        (terminated)
		.m_src_axi_rresp        (2'b00),                                                                //        (terminated)
		.m_src_axi_rdata        (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.m_src_axi_rready       (),                                                                     //        (terminated)
		.m_src_axi_awlen        (),                                                                     //        (terminated)
		.m_src_axi_awsize       (),                                                                     //        (terminated)
		.m_src_axi_awburst      (),                                                                     //        (terminated)
		.m_src_axi_awcache      (),                                                                     //        (terminated)
		.m_src_axi_awprot       (),                                                                     //        (terminated)
		.m_src_axi_wlast        (),                                                                     //        (terminated)
		.m_src_axi_arlen        (),                                                                     //        (terminated)
		.m_src_axi_arsize       (),                                                                     //        (terminated)
		.m_src_axi_arburst      (),                                                                     //        (terminated)
		.m_src_axi_arcache      (),                                                                     //        (terminated)
		.m_src_axi_arprot       (),                                                                     //        (terminated)
		.m_src_axi_awid         (),                                                                     //        (terminated)
		.m_src_axi_awlock       (),                                                                     //        (terminated)
		.m_src_axi_wid          (),                                                                     //        (terminated)
		.m_src_axi_arid         (),                                                                     //        (terminated)
		.m_src_axi_arlock       (),                                                                     //        (terminated)
		.m_src_axi_rid          (1'b0),                                                                 //        (terminated)
		.m_src_axi_bid          (1'b0),                                                                 //        (terminated)
		.m_src_axi_rlast        (1'b0)                                                                  //        (terminated)
	);

	spi_engine_execution #(
		.NUM_OF_CS       (1),
		.DEFAULT_SPI_CFG (0),
		.DEFAULT_CLK_DIV (0),
		.DATA_WIDTH      (18),
		.NUM_OF_SDI      (2),
		.SDO_DEFAULT     (2'b00),
		.SDI_DELAY       (3'b010)
	) spi_engine_execution_0 (
		.clk            (spi_engine_pll_outclk0_clk),                      //    clk.clk
		.resetn         (axi_spi_engine_0_spi_resetn_reset),               // resetn.reset_n
		.cmd_valid      (spi_engine_interconnect_0_m_ctrl_cmd_valid),      //   ctrl.cmd_valid
		.sdo_data_valid (spi_engine_interconnect_0_m_ctrl_sdo_data_valid), //       .sdo_data_valid
		.sdo_data_ready (spi_engine_execution_0_ctrl_sdo_data_ready),      //       .sdo_data_ready
		.sdo_data       (spi_engine_interconnect_0_m_ctrl_sdo_data),       //       .sdo_data
		.sdi_data_ready (spi_engine_interconnect_0_m_ctrl_sdi_data_ready), //       .sdi_data_ready
		.sdi_data_valid (spi_engine_execution_0_ctrl_sdi_data_valid),      //       .sdi_data_valid
		.sdi_data       (spi_engine_execution_0_ctrl_sdi_data),            //       .sdi_data
		.sync_ready     (spi_engine_interconnect_0_m_ctrl_sync_ready),     //       .sync_ready
		.sync_valid     (spi_engine_execution_0_ctrl_sync_valid),          //       .sync_valid
		.sync           (spi_engine_execution_0_ctrl_sync),                //       .sync
		.cmd_ready      (spi_engine_execution_0_ctrl_cmd_ready),           //       .cmd_ready
		.cmd            (spi_engine_interconnect_0_m_ctrl_cmd),            //       .cmd
		.three_wire     (spi_engine_execution_0_spi_out_three_wire),       //    spi.three_wire
		.sdo_t          (spi_engine_execution_0_spi_out_sdo_t),            //       .sdo_t
		.sdo            (spi_engine_execution_0_spi_out_sdo),              //       .sdo
		.sdi            (spi_engine_execution_0_spi_out_sdi),              //       .sdi
		.cs             (spi_engine_execution_0_spi_out_cs),               //       .cs
		.sclk           (spi_engine_execution_0_spi_out_sclk),             //       .sclk
		.sdi_1          (spi_engine_execution_0_spi_out_sdi_1),            //       .sdi_1
		.active         ()                                                 // active.active
	);

	spi_engine_interconnect #(
		.DATA_WIDTH (18),
		.NUM_OF_SDI (2)
	) spi_engine_interconnect_0 (
		.clk           (spi_engine_pll_outclk0_clk),                      //     clk.clk
		.resetn        (axi_spi_engine_0_spi_resetn_reset),               //  resetn.reset_n
		.s0_cmd_data   (spi_engine_offload_0_spi_engine_ctrl_cmd_data),   // s0_ctrl.cmd_data
		.s0_cmd_ready  (spi_engine_interconnect_0_s0_ctrl_cmd_ready),     //        .cmd_ready
		.s0_cmd_valid  (spi_engine_offload_0_spi_engine_ctrl_cmd_valid),  //        .cmd_valid
		.s0_sdo_data   (spi_engine_offload_0_spi_engine_ctrl_sdo_data),   //        .sdo_data
		.s0_sdo_valid  (spi_engine_offload_0_spi_engine_ctrl_sdo_valid),  //        .sdo_valid
		.s0_sdo_ready  (spi_engine_interconnect_0_s0_ctrl_sdo_ready),     //        .sdo_ready
		.s0_sdi_data   (spi_engine_interconnect_0_s0_ctrl_sdi_data),      //        .sdi_data
		.s0_sdi_valid  (spi_engine_interconnect_0_s0_ctrl_sdi_valid),     //        .sdi_valid
		.s0_sdi_ready  (spi_engine_offload_0_spi_engine_ctrl_sdi_ready),  //        .sdi_ready
		.s0_sync_ready (spi_engine_offload_0_spi_engine_ctrl_sync_ready), //        .sync_ready
		.s0_sync_valid (spi_engine_interconnect_0_s0_ctrl_sync_valid),    //        .sync_valid
		.s0_sync       (spi_engine_interconnect_0_s0_ctrl_sync_data),     //        .sync_data
		.s1_cmd_valid  (axi_spi_engine_0_spi_engine_ctrl_cmd_valid),      // s1_ctrl.cmd_valid
		.s1_cmd_ready  (spi_engine_interconnect_0_s1_ctrl_cmd_ready),     //        .cmd_ready
		.s1_cmd_data   (axi_spi_engine_0_spi_engine_ctrl_cmd_data),       //        .cmd_data
		.s1_sdo_valid  (axi_spi_engine_0_spi_engine_ctrl_sdo_valid),      //        .sdo_valid
		.s1_sdo_ready  (spi_engine_interconnect_0_s1_ctrl_sdo_ready),     //        .sdo_ready
		.s1_sdo_data   (axi_spi_engine_0_spi_engine_ctrl_sdo_data),       //        .sdo_data
		.s1_sdi_valid  (spi_engine_interconnect_0_s1_ctrl_sdi_valid),     //        .sdi_valid
		.s1_sdi_ready  (axi_spi_engine_0_spi_engine_ctrl_sdi_ready),      //        .sdi_ready
		.s1_sdi_data   (spi_engine_interconnect_0_s1_ctrl_sdi_data),      //        .sdi_data
		.s1_sync_valid (spi_engine_interconnect_0_s1_ctrl_sync_valid),    //        .sync_valid
		.s1_sync_ready (axi_spi_engine_0_spi_engine_ctrl_sync_ready),     //        .sync_ready
		.s1_sync       (spi_engine_interconnect_0_s1_ctrl_sync_data),     //        .sync_data
		.m_cmd_data    (spi_engine_interconnect_0_m_ctrl_cmd),            //  m_ctrl.cmd
		.m_cmd_valid   (spi_engine_interconnect_0_m_ctrl_cmd_valid),      //        .cmd_valid
		.m_cmd_ready   (spi_engine_execution_0_ctrl_cmd_ready),           //        .cmd_ready
		.m_sdo_valid   (spi_engine_interconnect_0_m_ctrl_sdo_data_valid), //        .sdo_data_valid
		.m_sdi_data    (spi_engine_execution_0_ctrl_sdi_data),            //        .sdi_data
		.m_sdi_valid   (spi_engine_execution_0_ctrl_sdi_data_valid),      //        .sdi_data_valid
		.m_sdi_ready   (spi_engine_interconnect_0_m_ctrl_sdi_data_ready), //        .sdi_data_ready
		.m_sdo_data    (spi_engine_interconnect_0_m_ctrl_sdo_data),       //        .sdo_data
		.m_sdo_ready   (spi_engine_execution_0_ctrl_sdo_data_ready),      //        .sdo_data_ready
		.m_sync        (spi_engine_execution_0_ctrl_sync),                //        .sync
		.m_sync_ready  (spi_engine_interconnect_0_m_ctrl_sync_ready),     //        .sync_ready
		.m_sync_valid  (spi_engine_execution_0_ctrl_sync_valid)           //        .sync_valid
	);

	spi_engine_offload #(
		.ASYNC_SPI_CLK         (1),
		.ASYNC_TRIG            (1),
		.CMD_MEM_ADDRESS_WIDTH (4),
		.SDO_MEM_ADDRESS_WIDTH (4),
		.DATA_WIDTH            (18),
		.NUM_OF_SDI            (2)
	) spi_engine_offload_0 (
		.ctrl_cmd_wr_en    (axi_spi_engine_0_spi_engine_offload_ctrl0_cmd_wr_en),   // spi_engine_offload_ctrl.cmd_wr_en
		.ctrl_cmd_wr_data  (axi_spi_engine_0_spi_engine_offload_ctrl0_cmd_wr_data), //                        .cmd_wr_data
		.ctrl_sdo_wr_en    (axi_spi_engine_0_spi_engine_offload_ctrl0_sdo_wr_en),   //                        .sdo_wr_en
		.ctrl_sdo_wr_data  (axi_spi_engine_0_spi_engine_offload_ctrl0_sdo_wr_data), //                        .sdo_wr_data
		.ctrl_enable       (axi_spi_engine_0_spi_engine_offload_ctrl0_enable),      //                        .enable
		.ctrl_enabled      (spi_engine_offload_0_spi_engine_offload_ctrl_enabled),  //                        .enabled
		.ctrl_mem_reset    (axi_spi_engine_0_spi_engine_offload_ctrl0_reset),       //                        .reset
		.ctrl_clk          (spi_engine_pll_outclk0_clk),                            //                ctrl_clk.clk
		.spi_clk           (spi_engine_pll_outclk0_clk),                            //                 spi_clk.clk
		.spi_resetn        (axi_spi_engine_0_spi_resetn_reset),                     //              spi_resetn.reset_n
		.trigger           (trigger_gen_0_pulse_pulse),                             //                 trigger.pulse
		.cmd_ready         (spi_engine_interconnect_0_s0_ctrl_cmd_ready),           //         spi_engine_ctrl.cmd_ready
		.cmd_valid         (spi_engine_offload_0_spi_engine_ctrl_cmd_valid),        //                        .cmd_valid
		.cmd               (spi_engine_offload_0_spi_engine_ctrl_cmd_data),         //                        .cmd_data
		.sdo_data_ready    (spi_engine_interconnect_0_s0_ctrl_sdo_ready),           //                        .sdo_ready
		.sdo_data_valid    (spi_engine_offload_0_spi_engine_ctrl_sdo_valid),        //                        .sdo_valid
		.sdo_data          (spi_engine_offload_0_spi_engine_ctrl_sdo_data),         //                        .sdo_data
		.sdi_data_ready    (spi_engine_offload_0_spi_engine_ctrl_sdi_ready),        //                        .sdi_ready
		.sdi_data_valid    (spi_engine_interconnect_0_s0_ctrl_sdi_valid),           //                        .sdi_valid
		.sdi_data          (spi_engine_interconnect_0_s0_ctrl_sdi_data),            //                        .sdi_data
		.sync_ready        (spi_engine_offload_0_spi_engine_ctrl_sync_ready),       //                        .sync_ready
		.sync_valid        (spi_engine_interconnect_0_s0_ctrl_sync_valid),          //                        .sync_valid
		.sync_data         (spi_engine_interconnect_0_s0_ctrl_sync_data),           //                        .sync_data
		.offload_sdi_ready (upscale_converter_0_s_axis_ready),                      //             offload_sdi.ready
		.offload_sdi_valid (spi_engine_offload_0_offload_sdi_valid),                //                        .valid
		.offload_sdi_data  (spi_engine_offload_0_offload_sdi_data)                  //                        .data
	);

	system_bd_spi_engine_pll spi_engine_pll (
		.refclk   (sys_hps_h2f_user1_clock_clk), //  refclk.clk
		.rst      (~sys_rst_reset_n),            //   reset.reset
		.outclk_0 (spi_engine_pll_outclk0_clk),  // outclk0.clk
		.locked   ()                             //  locked.export
	);

	system_bd_sys_gpio_bd sys_gpio_bd (
		.clk        (sys_hps_h2f_user1_clock_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_bd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_bd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_bd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_bd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_bd_s1_readdata),   //                    .readdata
		.in_port    (sys_gpio_bd_in_port),                         // external_connection.export
		.out_port   (sys_gpio_bd_out_port),                        //                    .export
		.irq        (irq_mapper_receiver2_irq)                     //                 irq.irq
	);

	system_bd_sys_gpio_in sys_gpio_in (
		.clk        (sys_hps_h2f_user1_clock_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_in_s1_readdata),   //                    .readdata
		.in_port    (sys_gpio_in_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                     //                 irq.irq
	);

	system_bd_sys_gpio_out sys_gpio_out (
		.clk        (sys_hps_h2f_user1_clock_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_out_s1_readdata),   //                    .readdata
		.out_port   (sys_gpio_out_export)                           // external_connection.export
	);

	system_bd_sys_hps #(
		.F2S_Width (2),
		.S2F_Width (2)
	) sys_hps (
		.h2f_user1_clk            (sys_hps_h2f_user1_clock_clk),                             //   h2f_user1_clock.clk
		.mem_a                    (sys_hps_memory_mem_a),                                    //            memory.mem_a
		.mem_ba                   (sys_hps_memory_mem_ba),                                   //                  .mem_ba
		.mem_ck                   (sys_hps_memory_mem_ck),                                   //                  .mem_ck
		.mem_ck_n                 (sys_hps_memory_mem_ck_n),                                 //                  .mem_ck_n
		.mem_cke                  (sys_hps_memory_mem_cke),                                  //                  .mem_cke
		.mem_cs_n                 (sys_hps_memory_mem_cs_n),                                 //                  .mem_cs_n
		.mem_ras_n                (sys_hps_memory_mem_ras_n),                                //                  .mem_ras_n
		.mem_cas_n                (sys_hps_memory_mem_cas_n),                                //                  .mem_cas_n
		.mem_we_n                 (sys_hps_memory_mem_we_n),                                 //                  .mem_we_n
		.mem_reset_n              (sys_hps_memory_mem_reset_n),                              //                  .mem_reset_n
		.mem_dq                   (sys_hps_memory_mem_dq),                                   //                  .mem_dq
		.mem_dqs                  (sys_hps_memory_mem_dqs),                                  //                  .mem_dqs
		.mem_dqs_n                (sys_hps_memory_mem_dqs_n),                                //                  .mem_dqs_n
		.mem_odt                  (sys_hps_memory_mem_odt),                                  //                  .mem_odt
		.mem_dm                   (sys_hps_memory_mem_dm),                                   //                  .mem_dm
		.oct_rzqin                (sys_hps_memory_oct_rzqin),                                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (sys_hps_hps_io_hps_io_emac1_inst_TX_CLK),                 //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (sys_hps_hps_io_hps_io_emac1_inst_TXD0),                   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (sys_hps_hps_io_hps_io_emac1_inst_TXD1),                   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (sys_hps_hps_io_hps_io_emac1_inst_TXD2),                   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (sys_hps_hps_io_hps_io_emac1_inst_TXD3),                   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (sys_hps_hps_io_hps_io_emac1_inst_RXD0),                   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (sys_hps_hps_io_hps_io_emac1_inst_MDIO),                   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (sys_hps_hps_io_hps_io_emac1_inst_MDC),                    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (sys_hps_hps_io_hps_io_emac1_inst_RX_CTL),                 //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (sys_hps_hps_io_hps_io_emac1_inst_TX_CTL),                 //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (sys_hps_hps_io_hps_io_emac1_inst_RX_CLK),                 //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (sys_hps_hps_io_hps_io_emac1_inst_RXD1),                   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (sys_hps_hps_io_hps_io_emac1_inst_RXD2),                   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (sys_hps_hps_io_hps_io_emac1_inst_RXD3),                   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (sys_hps_hps_io_hps_io_qspi_inst_IO0),                     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (sys_hps_hps_io_hps_io_qspi_inst_IO1),                     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (sys_hps_hps_io_hps_io_qspi_inst_IO2),                     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (sys_hps_hps_io_hps_io_qspi_inst_IO3),                     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (sys_hps_hps_io_hps_io_qspi_inst_SS0),                     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (sys_hps_hps_io_hps_io_qspi_inst_CLK),                     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (sys_hps_hps_io_hps_io_sdio_inst_CMD),                     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (sys_hps_hps_io_hps_io_sdio_inst_D0),                      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (sys_hps_hps_io_hps_io_sdio_inst_D1),                      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (sys_hps_hps_io_hps_io_sdio_inst_CLK),                     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (sys_hps_hps_io_hps_io_sdio_inst_D2),                      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (sys_hps_hps_io_hps_io_sdio_inst_D3),                      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (sys_hps_hps_io_hps_io_usb1_inst_D0),                      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (sys_hps_hps_io_hps_io_usb1_inst_D1),                      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (sys_hps_hps_io_hps_io_usb1_inst_D2),                      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (sys_hps_hps_io_hps_io_usb1_inst_D3),                      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (sys_hps_hps_io_hps_io_usb1_inst_D4),                      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (sys_hps_hps_io_hps_io_usb1_inst_D5),                      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (sys_hps_hps_io_hps_io_usb1_inst_D6),                      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (sys_hps_hps_io_hps_io_usb1_inst_D7),                      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (sys_hps_hps_io_hps_io_usb1_inst_CLK),                     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (sys_hps_hps_io_hps_io_usb1_inst_STP),                     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (sys_hps_hps_io_hps_io_usb1_inst_DIR),                     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (sys_hps_hps_io_hps_io_usb1_inst_NXT),                     //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (sys_hps_hps_io_hps_io_uart0_inst_RX),                     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (sys_hps_hps_io_hps_io_uart0_inst_TX),                     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (sys_hps_hps_io_hps_io_i2c0_inst_SDA),                     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (sys_hps_hps_io_hps_io_i2c0_inst_SCL),                     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (sys_hps_hps_io_hps_io_i2c1_inst_SDA),                     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (sys_hps_hps_io_hps_io_i2c1_inst_SCL),                     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO00  (sys_hps_hps_io_hps_io_gpio_inst_GPIO00),                  //                  .hps_io_gpio_inst_GPIO00
		.hps_io_gpio_inst_GPIO09  (sys_hps_hps_io_hps_io_gpio_inst_GPIO09),                  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (sys_hps_hps_io_hps_io_gpio_inst_GPIO35),                  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (sys_hps_hps_io_hps_io_gpio_inst_GPIO40),                  //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (sys_hps_hps_io_hps_io_gpio_inst_GPIO41),                  //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO42  (sys_hps_hps_io_hps_io_gpio_inst_GPIO42),                  //                  .hps_io_gpio_inst_GPIO42
		.hps_io_gpio_inst_GPIO43  (sys_hps_hps_io_hps_io_gpio_inst_GPIO43),                  //                  .hps_io_gpio_inst_GPIO43
		.hps_io_gpio_inst_GPIO44  (sys_hps_hps_io_hps_io_gpio_inst_GPIO44),                  //                  .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48  (sys_hps_hps_io_hps_io_gpio_inst_GPIO48),                  //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (sys_hps_hps_io_hps_io_gpio_inst_GPIO53),                  //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (sys_hps_hps_io_hps_io_gpio_inst_GPIO54),                  //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO55  (sys_hps_hps_io_hps_io_gpio_inst_GPIO55),                  //                  .hps_io_gpio_inst_GPIO55
		.hps_io_gpio_inst_GPIO56  (sys_hps_hps_io_hps_io_gpio_inst_GPIO56),                  //                  .hps_io_gpio_inst_GPIO56
		.hps_io_gpio_inst_GPIO57  (sys_hps_hps_io_hps_io_gpio_inst_GPIO57),                  //                  .hps_io_gpio_inst_GPIO57
		.hps_io_gpio_inst_GPIO58  (sys_hps_hps_io_hps_io_gpio_inst_GPIO58),                  //                  .hps_io_gpio_inst_GPIO58
		.hps_io_gpio_inst_GPIO59  (sys_hps_hps_io_hps_io_gpio_inst_GPIO59),                  //                  .hps_io_gpio_inst_GPIO59
		.hps_io_gpio_inst_GPIO61  (sys_hps_hps_io_hps_io_gpio_inst_GPIO61),                  //                  .hps_io_gpio_inst_GPIO61
		.hps_io_gpio_inst_GPIO65  (sys_hps_hps_io_hps_io_gpio_inst_GPIO65),                  //                  .hps_io_gpio_inst_GPIO65
		.h2f_rst_n                (sys_hps_h2f_reset_reset_n),                               //         h2f_reset.reset_n
		.f2h_sdram0_clk           (sys_hps_h2f_user1_clock_clk),                             //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_2_sys_hps_f2h_sdram0_data_address),       //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_2_sys_hps_f2h_sdram0_data_burstcount),    //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_2_sys_hps_f2h_sdram0_data_waitrequest),   //                  .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_2_sys_hps_f2h_sdram0_data_readdata),      //                  .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_2_sys_hps_f2h_sdram0_data_readdatavalid), //                  .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_2_sys_hps_f2h_sdram0_data_read),          //                  .read
		.f2h_sdram0_WRITEDATA     (mm_interconnect_2_sys_hps_f2h_sdram0_data_writedata),     //                  .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_2_sys_hps_f2h_sdram0_data_byteenable),    //                  .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_2_sys_hps_f2h_sdram0_data_write),         //                  .write
		.f2h_sdram1_clk           (sys_hps_h2f_user1_clock_clk),                             //  f2h_sdram1_clock.clk
		.f2h_sdram1_ARADDR        (mm_interconnect_1_sys_hps_f2h_sdram1_data_araddr),        //   f2h_sdram1_data.araddr
		.f2h_sdram1_ARLEN         (mm_interconnect_1_sys_hps_f2h_sdram1_data_arlen),         //                  .arlen
		.f2h_sdram1_ARID          (mm_interconnect_1_sys_hps_f2h_sdram1_data_arid),          //                  .arid
		.f2h_sdram1_ARSIZE        (mm_interconnect_1_sys_hps_f2h_sdram1_data_arsize),        //                  .arsize
		.f2h_sdram1_ARBURST       (mm_interconnect_1_sys_hps_f2h_sdram1_data_arburst),       //                  .arburst
		.f2h_sdram1_ARLOCK        (mm_interconnect_1_sys_hps_f2h_sdram1_data_arlock),        //                  .arlock
		.f2h_sdram1_ARPROT        (mm_interconnect_1_sys_hps_f2h_sdram1_data_arprot),        //                  .arprot
		.f2h_sdram1_ARVALID       (mm_interconnect_1_sys_hps_f2h_sdram1_data_arvalid),       //                  .arvalid
		.f2h_sdram1_ARCACHE       (mm_interconnect_1_sys_hps_f2h_sdram1_data_arcache),       //                  .arcache
		.f2h_sdram1_AWADDR        (mm_interconnect_1_sys_hps_f2h_sdram1_data_awaddr),        //                  .awaddr
		.f2h_sdram1_AWLEN         (mm_interconnect_1_sys_hps_f2h_sdram1_data_awlen),         //                  .awlen
		.f2h_sdram1_AWID          (mm_interconnect_1_sys_hps_f2h_sdram1_data_awid),          //                  .awid
		.f2h_sdram1_AWSIZE        (mm_interconnect_1_sys_hps_f2h_sdram1_data_awsize),        //                  .awsize
		.f2h_sdram1_AWBURST       (mm_interconnect_1_sys_hps_f2h_sdram1_data_awburst),       //                  .awburst
		.f2h_sdram1_AWLOCK        (mm_interconnect_1_sys_hps_f2h_sdram1_data_awlock),        //                  .awlock
		.f2h_sdram1_AWPROT        (mm_interconnect_1_sys_hps_f2h_sdram1_data_awprot),        //                  .awprot
		.f2h_sdram1_AWVALID       (mm_interconnect_1_sys_hps_f2h_sdram1_data_awvalid),       //                  .awvalid
		.f2h_sdram1_AWCACHE       (mm_interconnect_1_sys_hps_f2h_sdram1_data_awcache),       //                  .awcache
		.f2h_sdram1_BRESP         (mm_interconnect_1_sys_hps_f2h_sdram1_data_bresp),         //                  .bresp
		.f2h_sdram1_BID           (mm_interconnect_1_sys_hps_f2h_sdram1_data_bid),           //                  .bid
		.f2h_sdram1_BVALID        (mm_interconnect_1_sys_hps_f2h_sdram1_data_bvalid),        //                  .bvalid
		.f2h_sdram1_BREADY        (mm_interconnect_1_sys_hps_f2h_sdram1_data_bready),        //                  .bready
		.f2h_sdram1_ARREADY       (mm_interconnect_1_sys_hps_f2h_sdram1_data_arready),       //                  .arready
		.f2h_sdram1_AWREADY       (mm_interconnect_1_sys_hps_f2h_sdram1_data_awready),       //                  .awready
		.f2h_sdram1_RREADY        (mm_interconnect_1_sys_hps_f2h_sdram1_data_rready),        //                  .rready
		.f2h_sdram1_RDATA         (mm_interconnect_1_sys_hps_f2h_sdram1_data_rdata),         //                  .rdata
		.f2h_sdram1_RRESP         (mm_interconnect_1_sys_hps_f2h_sdram1_data_rresp),         //                  .rresp
		.f2h_sdram1_RLAST         (mm_interconnect_1_sys_hps_f2h_sdram1_data_rlast),         //                  .rlast
		.f2h_sdram1_RID           (mm_interconnect_1_sys_hps_f2h_sdram1_data_rid),           //                  .rid
		.f2h_sdram1_RVALID        (mm_interconnect_1_sys_hps_f2h_sdram1_data_rvalid),        //                  .rvalid
		.f2h_sdram1_WLAST         (mm_interconnect_1_sys_hps_f2h_sdram1_data_wlast),         //                  .wlast
		.f2h_sdram1_WVALID        (mm_interconnect_1_sys_hps_f2h_sdram1_data_wvalid),        //                  .wvalid
		.f2h_sdram1_WDATA         (mm_interconnect_1_sys_hps_f2h_sdram1_data_wdata),         //                  .wdata
		.f2h_sdram1_WSTRB         (mm_interconnect_1_sys_hps_f2h_sdram1_data_wstrb),         //                  .wstrb
		.f2h_sdram1_WREADY        (mm_interconnect_1_sys_hps_f2h_sdram1_data_wready),        //                  .wready
		.f2h_sdram1_WID           (mm_interconnect_1_sys_hps_f2h_sdram1_data_wid),           //                  .wid
		.f2h_sdram2_clk           (sys_hps_h2f_user1_clock_clk),                             //  f2h_sdram2_clock.clk
		.f2h_sdram2_ARADDR        (),                                                        //   f2h_sdram2_data.araddr
		.f2h_sdram2_ARLEN         (),                                                        //                  .arlen
		.f2h_sdram2_ARID          (),                                                        //                  .arid
		.f2h_sdram2_ARSIZE        (),                                                        //                  .arsize
		.f2h_sdram2_ARBURST       (),                                                        //                  .arburst
		.f2h_sdram2_ARLOCK        (),                                                        //                  .arlock
		.f2h_sdram2_ARPROT        (),                                                        //                  .arprot
		.f2h_sdram2_ARVALID       (),                                                        //                  .arvalid
		.f2h_sdram2_ARCACHE       (),                                                        //                  .arcache
		.f2h_sdram2_AWADDR        (),                                                        //                  .awaddr
		.f2h_sdram2_AWLEN         (),                                                        //                  .awlen
		.f2h_sdram2_AWID          (),                                                        //                  .awid
		.f2h_sdram2_AWSIZE        (),                                                        //                  .awsize
		.f2h_sdram2_AWBURST       (),                                                        //                  .awburst
		.f2h_sdram2_AWLOCK        (),                                                        //                  .awlock
		.f2h_sdram2_AWPROT        (),                                                        //                  .awprot
		.f2h_sdram2_AWVALID       (),                                                        //                  .awvalid
		.f2h_sdram2_AWCACHE       (),                                                        //                  .awcache
		.f2h_sdram2_BRESP         (),                                                        //                  .bresp
		.f2h_sdram2_BID           (),                                                        //                  .bid
		.f2h_sdram2_BVALID        (),                                                        //                  .bvalid
		.f2h_sdram2_BREADY        (),                                                        //                  .bready
		.f2h_sdram2_ARREADY       (),                                                        //                  .arready
		.f2h_sdram2_AWREADY       (),                                                        //                  .awready
		.f2h_sdram2_RREADY        (),                                                        //                  .rready
		.f2h_sdram2_RDATA         (),                                                        //                  .rdata
		.f2h_sdram2_RRESP         (),                                                        //                  .rresp
		.f2h_sdram2_RLAST         (),                                                        //                  .rlast
		.f2h_sdram2_RID           (),                                                        //                  .rid
		.f2h_sdram2_RVALID        (),                                                        //                  .rvalid
		.f2h_sdram2_WLAST         (),                                                        //                  .wlast
		.f2h_sdram2_WVALID        (),                                                        //                  .wvalid
		.f2h_sdram2_WDATA         (),                                                        //                  .wdata
		.f2h_sdram2_WSTRB         (),                                                        //                  .wstrb
		.f2h_sdram2_WREADY        (),                                                        //                  .wready
		.f2h_sdram2_WID           (),                                                        //                  .wid
		.h2f_axi_clk              (sys_hps_h2f_user1_clock_clk),                             //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                                        //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                                        //                  .awaddr
		.h2f_AWLEN                (),                                                        //                  .awlen
		.h2f_AWSIZE               (),                                                        //                  .awsize
		.h2f_AWBURST              (),                                                        //                  .awburst
		.h2f_AWLOCK               (),                                                        //                  .awlock
		.h2f_AWCACHE              (),                                                        //                  .awcache
		.h2f_AWPROT               (),                                                        //                  .awprot
		.h2f_AWVALID              (),                                                        //                  .awvalid
		.h2f_AWREADY              (),                                                        //                  .awready
		.h2f_WID                  (),                                                        //                  .wid
		.h2f_WDATA                (),                                                        //                  .wdata
		.h2f_WSTRB                (),                                                        //                  .wstrb
		.h2f_WLAST                (),                                                        //                  .wlast
		.h2f_WVALID               (),                                                        //                  .wvalid
		.h2f_WREADY               (),                                                        //                  .wready
		.h2f_BID                  (),                                                        //                  .bid
		.h2f_BRESP                (),                                                        //                  .bresp
		.h2f_BVALID               (),                                                        //                  .bvalid
		.h2f_BREADY               (),                                                        //                  .bready
		.h2f_ARID                 (),                                                        //                  .arid
		.h2f_ARADDR               (),                                                        //                  .araddr
		.h2f_ARLEN                (),                                                        //                  .arlen
		.h2f_ARSIZE               (),                                                        //                  .arsize
		.h2f_ARBURST              (),                                                        //                  .arburst
		.h2f_ARLOCK               (),                                                        //                  .arlock
		.h2f_ARCACHE              (),                                                        //                  .arcache
		.h2f_ARPROT               (),                                                        //                  .arprot
		.h2f_ARVALID              (),                                                        //                  .arvalid
		.h2f_ARREADY              (),                                                        //                  .arready
		.h2f_RID                  (),                                                        //                  .rid
		.h2f_RDATA                (),                                                        //                  .rdata
		.h2f_RRESP                (),                                                        //                  .rresp
		.h2f_RLAST                (),                                                        //                  .rlast
		.h2f_RVALID               (),                                                        //                  .rvalid
		.h2f_RREADY               (),                                                        //                  .rready
		.f2h_axi_clk              (sys_hps_h2f_user1_clock_clk),                             //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                                        //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                                        //                  .awaddr
		.f2h_AWLEN                (),                                                        //                  .awlen
		.f2h_AWSIZE               (),                                                        //                  .awsize
		.f2h_AWBURST              (),                                                        //                  .awburst
		.f2h_AWLOCK               (),                                                        //                  .awlock
		.f2h_AWCACHE              (),                                                        //                  .awcache
		.f2h_AWPROT               (),                                                        //                  .awprot
		.f2h_AWVALID              (),                                                        //                  .awvalid
		.f2h_AWREADY              (),                                                        //                  .awready
		.f2h_AWUSER               (),                                                        //                  .awuser
		.f2h_WID                  (),                                                        //                  .wid
		.f2h_WDATA                (),                                                        //                  .wdata
		.f2h_WSTRB                (),                                                        //                  .wstrb
		.f2h_WLAST                (),                                                        //                  .wlast
		.f2h_WVALID               (),                                                        //                  .wvalid
		.f2h_WREADY               (),                                                        //                  .wready
		.f2h_BID                  (),                                                        //                  .bid
		.f2h_BRESP                (),                                                        //                  .bresp
		.f2h_BVALID               (),                                                        //                  .bvalid
		.f2h_BREADY               (),                                                        //                  .bready
		.f2h_ARID                 (),                                                        //                  .arid
		.f2h_ARADDR               (),                                                        //                  .araddr
		.f2h_ARLEN                (),                                                        //                  .arlen
		.f2h_ARSIZE               (),                                                        //                  .arsize
		.f2h_ARBURST              (),                                                        //                  .arburst
		.f2h_ARLOCK               (),                                                        //                  .arlock
		.f2h_ARCACHE              (),                                                        //                  .arcache
		.f2h_ARPROT               (),                                                        //                  .arprot
		.f2h_ARVALID              (),                                                        //                  .arvalid
		.f2h_ARREADY              (),                                                        //                  .arready
		.f2h_ARUSER               (),                                                        //                  .aruser
		.f2h_RID                  (),                                                        //                  .rid
		.f2h_RDATA                (),                                                        //                  .rdata
		.f2h_RRESP                (),                                                        //                  .rresp
		.f2h_RLAST                (),                                                        //                  .rlast
		.f2h_RVALID               (),                                                        //                  .rvalid
		.f2h_RREADY               (),                                                        //                  .rready
		.h2f_lw_axi_clk           (sys_hps_h2f_user1_clock_clk),                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (sys_hps_h2f_lw_axi_master_awid),                          // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (sys_hps_h2f_lw_axi_master_awaddr),                        //                  .awaddr
		.h2f_lw_AWLEN             (sys_hps_h2f_lw_axi_master_awlen),                         //                  .awlen
		.h2f_lw_AWSIZE            (sys_hps_h2f_lw_axi_master_awsize),                        //                  .awsize
		.h2f_lw_AWBURST           (sys_hps_h2f_lw_axi_master_awburst),                       //                  .awburst
		.h2f_lw_AWLOCK            (sys_hps_h2f_lw_axi_master_awlock),                        //                  .awlock
		.h2f_lw_AWCACHE           (sys_hps_h2f_lw_axi_master_awcache),                       //                  .awcache
		.h2f_lw_AWPROT            (sys_hps_h2f_lw_axi_master_awprot),                        //                  .awprot
		.h2f_lw_AWVALID           (sys_hps_h2f_lw_axi_master_awvalid),                       //                  .awvalid
		.h2f_lw_AWREADY           (sys_hps_h2f_lw_axi_master_awready),                       //                  .awready
		.h2f_lw_WID               (sys_hps_h2f_lw_axi_master_wid),                           //                  .wid
		.h2f_lw_WDATA             (sys_hps_h2f_lw_axi_master_wdata),                         //                  .wdata
		.h2f_lw_WSTRB             (sys_hps_h2f_lw_axi_master_wstrb),                         //                  .wstrb
		.h2f_lw_WLAST             (sys_hps_h2f_lw_axi_master_wlast),                         //                  .wlast
		.h2f_lw_WVALID            (sys_hps_h2f_lw_axi_master_wvalid),                        //                  .wvalid
		.h2f_lw_WREADY            (sys_hps_h2f_lw_axi_master_wready),                        //                  .wready
		.h2f_lw_BID               (sys_hps_h2f_lw_axi_master_bid),                           //                  .bid
		.h2f_lw_BRESP             (sys_hps_h2f_lw_axi_master_bresp),                         //                  .bresp
		.h2f_lw_BVALID            (sys_hps_h2f_lw_axi_master_bvalid),                        //                  .bvalid
		.h2f_lw_BREADY            (sys_hps_h2f_lw_axi_master_bready),                        //                  .bready
		.h2f_lw_ARID              (sys_hps_h2f_lw_axi_master_arid),                          //                  .arid
		.h2f_lw_ARADDR            (sys_hps_h2f_lw_axi_master_araddr),                        //                  .araddr
		.h2f_lw_ARLEN             (sys_hps_h2f_lw_axi_master_arlen),                         //                  .arlen
		.h2f_lw_ARSIZE            (sys_hps_h2f_lw_axi_master_arsize),                        //                  .arsize
		.h2f_lw_ARBURST           (sys_hps_h2f_lw_axi_master_arburst),                       //                  .arburst
		.h2f_lw_ARLOCK            (sys_hps_h2f_lw_axi_master_arlock),                        //                  .arlock
		.h2f_lw_ARCACHE           (sys_hps_h2f_lw_axi_master_arcache),                       //                  .arcache
		.h2f_lw_ARPROT            (sys_hps_h2f_lw_axi_master_arprot),                        //                  .arprot
		.h2f_lw_ARVALID           (sys_hps_h2f_lw_axi_master_arvalid),                       //                  .arvalid
		.h2f_lw_ARREADY           (sys_hps_h2f_lw_axi_master_arready),                       //                  .arready
		.h2f_lw_RID               (sys_hps_h2f_lw_axi_master_rid),                           //                  .rid
		.h2f_lw_RDATA             (sys_hps_h2f_lw_axi_master_rdata),                         //                  .rdata
		.h2f_lw_RRESP             (sys_hps_h2f_lw_axi_master_rresp),                         //                  .rresp
		.h2f_lw_RLAST             (sys_hps_h2f_lw_axi_master_rlast),                         //                  .rlast
		.h2f_lw_RVALID            (sys_hps_h2f_lw_axi_master_rvalid),                        //                  .rvalid
		.h2f_lw_RREADY            (sys_hps_h2f_lw_axi_master_rready),                        //                  .rready
		.f2h_irq_p0               (sys_hps_f2h_irq0_irq),                                    //          f2h_irq0.irq
		.f2h_irq_p1               (sys_hps_f2h_irq1_irq)                                     //          f2h_irq1.irq
	);

	system_bd_sys_id sys_id (
		.clock    (sys_hps_h2f_user1_clock_clk),                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	util_pulse_gen #(
		.PULSE_PERIOD (40),
		.PULSE_WIDTH  (1)
	) trigger_gen_0 (
		.clk           (spi_engine_pll_outclk0_clk),              //           clk.clk
		.rstn          (axi_spi_engine_0_spi_resetn_reset),       //          rstn.reset_n
		.pulse_width   (trigger_gen_0_pulse_width_pulse_width),   //   pulse_width.pulse_width
		.pulse_period  (trigger_gen_0_pulse_period_pulse_period), //  pulse_period.pulse_period
		.load_config   (trigger_gen_0_load_config_load_config),   //   load_config.load_config
		.pulse         (trigger_gen_0_pulse_pulse),               //         pulse.pulse
		.pulse_counter ()                                         // pulse_counter.pulse_counter
	);

	util_axis_upscale_2 #(
		.NUM_OF_CHANNELS (2),
		.DATA_WIDTH      (18),
		.UDATA_WIDTH     (32)
	) upscale_converter_0 (
		.clk          (spi_engine_pll_outclk0_clk),                  //         clk.clk
		.resetn       (axi_spi_engine_0_spi_resetn_reset),           //      resetn.reset_n
		.dfmt_enable  (upscale_converter_0_dfmt_enable_dfmt_enable), // dfmt_enable.dfmt_enable
		.dfmt_se      (upscale_converter_0_dfmt_se_dfmt_se),         //     dfmt_se.dfmt_se
		.dfmt_type    (upscale_converter_0_dfmt_type_dfmt_type),     //   dfmt_type.dfmt_type
		.m_axis_data  (upscale_converter_0_m_axis_tdata),            //      m_axis.tdata
		.m_axis_ready (upscale_converter_0_m_axis_tready),           //            .tready
		.m_axis_valid (upscale_converter_0_m_axis_tvalid),           //            .tvalid
		.s_axis_valid (spi_engine_offload_0_offload_sdi_valid),      //      s_axis.valid
		.s_axis_ready (upscale_converter_0_s_axis_ready),            //            .ready
		.s_axis_data  (spi_engine_offload_0_offload_sdi_data)        //            .data
	);

	system_bd_mm_interconnect_0 mm_interconnect_0 (
		.axi_hdmi_tx_0_s_axi_awaddr                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awaddr),     //                                             axi_hdmi_tx_0_s_axi.awaddr
		.axi_hdmi_tx_0_s_axi_awprot                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awprot),     //                                                                .awprot
		.axi_hdmi_tx_0_s_axi_awvalid                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awvalid),    //                                                                .awvalid
		.axi_hdmi_tx_0_s_axi_awready                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awready),    //                                                                .awready
		.axi_hdmi_tx_0_s_axi_wdata                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wdata),      //                                                                .wdata
		.axi_hdmi_tx_0_s_axi_wstrb                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wstrb),      //                                                                .wstrb
		.axi_hdmi_tx_0_s_axi_wvalid                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wvalid),     //                                                                .wvalid
		.axi_hdmi_tx_0_s_axi_wready                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wready),     //                                                                .wready
		.axi_hdmi_tx_0_s_axi_bresp                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bresp),      //                                                                .bresp
		.axi_hdmi_tx_0_s_axi_bvalid                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bvalid),     //                                                                .bvalid
		.axi_hdmi_tx_0_s_axi_bready                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bready),     //                                                                .bready
		.axi_hdmi_tx_0_s_axi_araddr                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_araddr),     //                                                                .araddr
		.axi_hdmi_tx_0_s_axi_arprot                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arprot),     //                                                                .arprot
		.axi_hdmi_tx_0_s_axi_arvalid                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arvalid),    //                                                                .arvalid
		.axi_hdmi_tx_0_s_axi_arready                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arready),    //                                                                .arready
		.axi_hdmi_tx_0_s_axi_rdata                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rdata),      //                                                                .rdata
		.axi_hdmi_tx_0_s_axi_rresp                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rresp),      //                                                                .rresp
		.axi_hdmi_tx_0_s_axi_rvalid                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rvalid),     //                                                                .rvalid
		.axi_hdmi_tx_0_s_axi_rready                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rready),     //                                                                .rready
		.axi_spi_engine_0_s_axi_awaddr                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_awaddr),  //                                          axi_spi_engine_0_s_axi.awaddr
		.axi_spi_engine_0_s_axi_awprot                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_awprot),  //                                                                .awprot
		.axi_spi_engine_0_s_axi_awvalid                                        (mm_interconnect_0_axi_spi_engine_0_s_axi_awvalid), //                                                                .awvalid
		.axi_spi_engine_0_s_axi_awready                                        (mm_interconnect_0_axi_spi_engine_0_s_axi_awready), //                                                                .awready
		.axi_spi_engine_0_s_axi_wdata                                          (mm_interconnect_0_axi_spi_engine_0_s_axi_wdata),   //                                                                .wdata
		.axi_spi_engine_0_s_axi_wstrb                                          (mm_interconnect_0_axi_spi_engine_0_s_axi_wstrb),   //                                                                .wstrb
		.axi_spi_engine_0_s_axi_wvalid                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_wvalid),  //                                                                .wvalid
		.axi_spi_engine_0_s_axi_wready                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_wready),  //                                                                .wready
		.axi_spi_engine_0_s_axi_bresp                                          (mm_interconnect_0_axi_spi_engine_0_s_axi_bresp),   //                                                                .bresp
		.axi_spi_engine_0_s_axi_bvalid                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_bvalid),  //                                                                .bvalid
		.axi_spi_engine_0_s_axi_bready                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_bready),  //                                                                .bready
		.axi_spi_engine_0_s_axi_araddr                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_araddr),  //                                                                .araddr
		.axi_spi_engine_0_s_axi_arprot                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_arprot),  //                                                                .arprot
		.axi_spi_engine_0_s_axi_arvalid                                        (mm_interconnect_0_axi_spi_engine_0_s_axi_arvalid), //                                                                .arvalid
		.axi_spi_engine_0_s_axi_arready                                        (mm_interconnect_0_axi_spi_engine_0_s_axi_arready), //                                                                .arready
		.axi_spi_engine_0_s_axi_rdata                                          (mm_interconnect_0_axi_spi_engine_0_s_axi_rdata),   //                                                                .rdata
		.axi_spi_engine_0_s_axi_rresp                                          (mm_interconnect_0_axi_spi_engine_0_s_axi_rresp),   //                                                                .rresp
		.axi_spi_engine_0_s_axi_rvalid                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_rvalid),  //                                                                .rvalid
		.axi_spi_engine_0_s_axi_rready                                         (mm_interconnect_0_axi_spi_engine_0_s_axi_rready),  //                                                                .rready
		.hdmi_dmac_0_s_axi_awaddr                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_awaddr),       //                                               hdmi_dmac_0_s_axi.awaddr
		.hdmi_dmac_0_s_axi_awprot                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_awprot),       //                                                                .awprot
		.hdmi_dmac_0_s_axi_awvalid                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_awvalid),      //                                                                .awvalid
		.hdmi_dmac_0_s_axi_awready                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_awready),      //                                                                .awready
		.hdmi_dmac_0_s_axi_wdata                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_wdata),        //                                                                .wdata
		.hdmi_dmac_0_s_axi_wstrb                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_wstrb),        //                                                                .wstrb
		.hdmi_dmac_0_s_axi_wvalid                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_wvalid),       //                                                                .wvalid
		.hdmi_dmac_0_s_axi_wready                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_wready),       //                                                                .wready
		.hdmi_dmac_0_s_axi_bresp                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_bresp),        //                                                                .bresp
		.hdmi_dmac_0_s_axi_bvalid                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_bvalid),       //                                                                .bvalid
		.hdmi_dmac_0_s_axi_bready                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_bready),       //                                                                .bready
		.hdmi_dmac_0_s_axi_araddr                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_araddr),       //                                                                .araddr
		.hdmi_dmac_0_s_axi_arprot                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_arprot),       //                                                                .arprot
		.hdmi_dmac_0_s_axi_arvalid                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_arvalid),      //                                                                .arvalid
		.hdmi_dmac_0_s_axi_arready                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_arready),      //                                                                .arready
		.hdmi_dmac_0_s_axi_rdata                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_rdata),        //                                                                .rdata
		.hdmi_dmac_0_s_axi_rresp                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_rresp),        //                                                                .rresp
		.hdmi_dmac_0_s_axi_rvalid                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_rvalid),       //                                                                .rvalid
		.hdmi_dmac_0_s_axi_rready                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_rready),       //                                                                .rready
		.spi_dmac_0_s_axi_awaddr                                               (mm_interconnect_0_spi_dmac_0_s_axi_awaddr),        //                                                spi_dmac_0_s_axi.awaddr
		.spi_dmac_0_s_axi_awprot                                               (mm_interconnect_0_spi_dmac_0_s_axi_awprot),        //                                                                .awprot
		.spi_dmac_0_s_axi_awvalid                                              (mm_interconnect_0_spi_dmac_0_s_axi_awvalid),       //                                                                .awvalid
		.spi_dmac_0_s_axi_awready                                              (mm_interconnect_0_spi_dmac_0_s_axi_awready),       //                                                                .awready
		.spi_dmac_0_s_axi_wdata                                                (mm_interconnect_0_spi_dmac_0_s_axi_wdata),         //                                                                .wdata
		.spi_dmac_0_s_axi_wstrb                                                (mm_interconnect_0_spi_dmac_0_s_axi_wstrb),         //                                                                .wstrb
		.spi_dmac_0_s_axi_wvalid                                               (mm_interconnect_0_spi_dmac_0_s_axi_wvalid),        //                                                                .wvalid
		.spi_dmac_0_s_axi_wready                                               (mm_interconnect_0_spi_dmac_0_s_axi_wready),        //                                                                .wready
		.spi_dmac_0_s_axi_bresp                                                (mm_interconnect_0_spi_dmac_0_s_axi_bresp),         //                                                                .bresp
		.spi_dmac_0_s_axi_bvalid                                               (mm_interconnect_0_spi_dmac_0_s_axi_bvalid),        //                                                                .bvalid
		.spi_dmac_0_s_axi_bready                                               (mm_interconnect_0_spi_dmac_0_s_axi_bready),        //                                                                .bready
		.spi_dmac_0_s_axi_araddr                                               (mm_interconnect_0_spi_dmac_0_s_axi_araddr),        //                                                                .araddr
		.spi_dmac_0_s_axi_arprot                                               (mm_interconnect_0_spi_dmac_0_s_axi_arprot),        //                                                                .arprot
		.spi_dmac_0_s_axi_arvalid                                              (mm_interconnect_0_spi_dmac_0_s_axi_arvalid),       //                                                                .arvalid
		.spi_dmac_0_s_axi_arready                                              (mm_interconnect_0_spi_dmac_0_s_axi_arready),       //                                                                .arready
		.spi_dmac_0_s_axi_rdata                                                (mm_interconnect_0_spi_dmac_0_s_axi_rdata),         //                                                                .rdata
		.spi_dmac_0_s_axi_rresp                                                (mm_interconnect_0_spi_dmac_0_s_axi_rresp),         //                                                                .rresp
		.spi_dmac_0_s_axi_rvalid                                               (mm_interconnect_0_spi_dmac_0_s_axi_rvalid),        //                                                                .rvalid
		.spi_dmac_0_s_axi_rready                                               (mm_interconnect_0_spi_dmac_0_s_axi_rready),        //                                                                .rready
		.sys_hps_h2f_lw_axi_master_awid                                        (sys_hps_h2f_lw_axi_master_awid),                   //                                       sys_hps_h2f_lw_axi_master.awid
		.sys_hps_h2f_lw_axi_master_awaddr                                      (sys_hps_h2f_lw_axi_master_awaddr),                 //                                                                .awaddr
		.sys_hps_h2f_lw_axi_master_awlen                                       (sys_hps_h2f_lw_axi_master_awlen),                  //                                                                .awlen
		.sys_hps_h2f_lw_axi_master_awsize                                      (sys_hps_h2f_lw_axi_master_awsize),                 //                                                                .awsize
		.sys_hps_h2f_lw_axi_master_awburst                                     (sys_hps_h2f_lw_axi_master_awburst),                //                                                                .awburst
		.sys_hps_h2f_lw_axi_master_awlock                                      (sys_hps_h2f_lw_axi_master_awlock),                 //                                                                .awlock
		.sys_hps_h2f_lw_axi_master_awcache                                     (sys_hps_h2f_lw_axi_master_awcache),                //                                                                .awcache
		.sys_hps_h2f_lw_axi_master_awprot                                      (sys_hps_h2f_lw_axi_master_awprot),                 //                                                                .awprot
		.sys_hps_h2f_lw_axi_master_awvalid                                     (sys_hps_h2f_lw_axi_master_awvalid),                //                                                                .awvalid
		.sys_hps_h2f_lw_axi_master_awready                                     (sys_hps_h2f_lw_axi_master_awready),                //                                                                .awready
		.sys_hps_h2f_lw_axi_master_wid                                         (sys_hps_h2f_lw_axi_master_wid),                    //                                                                .wid
		.sys_hps_h2f_lw_axi_master_wdata                                       (sys_hps_h2f_lw_axi_master_wdata),                  //                                                                .wdata
		.sys_hps_h2f_lw_axi_master_wstrb                                       (sys_hps_h2f_lw_axi_master_wstrb),                  //                                                                .wstrb
		.sys_hps_h2f_lw_axi_master_wlast                                       (sys_hps_h2f_lw_axi_master_wlast),                  //                                                                .wlast
		.sys_hps_h2f_lw_axi_master_wvalid                                      (sys_hps_h2f_lw_axi_master_wvalid),                 //                                                                .wvalid
		.sys_hps_h2f_lw_axi_master_wready                                      (sys_hps_h2f_lw_axi_master_wready),                 //                                                                .wready
		.sys_hps_h2f_lw_axi_master_bid                                         (sys_hps_h2f_lw_axi_master_bid),                    //                                                                .bid
		.sys_hps_h2f_lw_axi_master_bresp                                       (sys_hps_h2f_lw_axi_master_bresp),                  //                                                                .bresp
		.sys_hps_h2f_lw_axi_master_bvalid                                      (sys_hps_h2f_lw_axi_master_bvalid),                 //                                                                .bvalid
		.sys_hps_h2f_lw_axi_master_bready                                      (sys_hps_h2f_lw_axi_master_bready),                 //                                                                .bready
		.sys_hps_h2f_lw_axi_master_arid                                        (sys_hps_h2f_lw_axi_master_arid),                   //                                                                .arid
		.sys_hps_h2f_lw_axi_master_araddr                                      (sys_hps_h2f_lw_axi_master_araddr),                 //                                                                .araddr
		.sys_hps_h2f_lw_axi_master_arlen                                       (sys_hps_h2f_lw_axi_master_arlen),                  //                                                                .arlen
		.sys_hps_h2f_lw_axi_master_arsize                                      (sys_hps_h2f_lw_axi_master_arsize),                 //                                                                .arsize
		.sys_hps_h2f_lw_axi_master_arburst                                     (sys_hps_h2f_lw_axi_master_arburst),                //                                                                .arburst
		.sys_hps_h2f_lw_axi_master_arlock                                      (sys_hps_h2f_lw_axi_master_arlock),                 //                                                                .arlock
		.sys_hps_h2f_lw_axi_master_arcache                                     (sys_hps_h2f_lw_axi_master_arcache),                //                                                                .arcache
		.sys_hps_h2f_lw_axi_master_arprot                                      (sys_hps_h2f_lw_axi_master_arprot),                 //                                                                .arprot
		.sys_hps_h2f_lw_axi_master_arvalid                                     (sys_hps_h2f_lw_axi_master_arvalid),                //                                                                .arvalid
		.sys_hps_h2f_lw_axi_master_arready                                     (sys_hps_h2f_lw_axi_master_arready),                //                                                                .arready
		.sys_hps_h2f_lw_axi_master_rid                                         (sys_hps_h2f_lw_axi_master_rid),                    //                                                                .rid
		.sys_hps_h2f_lw_axi_master_rdata                                       (sys_hps_h2f_lw_axi_master_rdata),                  //                                                                .rdata
		.sys_hps_h2f_lw_axi_master_rresp                                       (sys_hps_h2f_lw_axi_master_rresp),                  //                                                                .rresp
		.sys_hps_h2f_lw_axi_master_rlast                                       (sys_hps_h2f_lw_axi_master_rlast),                  //                                                                .rlast
		.sys_hps_h2f_lw_axi_master_rvalid                                      (sys_hps_h2f_lw_axi_master_rvalid),                 //                                                                .rvalid
		.sys_hps_h2f_lw_axi_master_rready                                      (sys_hps_h2f_lw_axi_master_rready),                 //                                                                .rready
		.sys_hps_h2f_user1_clock_clk                                           (sys_hps_h2f_user1_clock_clk),                      //                                         sys_hps_h2f_user1_clock.clk
		.sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),               // sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sys_id_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                   //                              sys_id_reset_reset_bridge_in_reset.reset
		.sys_gpio_bd_s1_address                                                (mm_interconnect_0_sys_gpio_bd_s1_address),         //                                                  sys_gpio_bd_s1.address
		.sys_gpio_bd_s1_write                                                  (mm_interconnect_0_sys_gpio_bd_s1_write),           //                                                                .write
		.sys_gpio_bd_s1_readdata                                               (mm_interconnect_0_sys_gpio_bd_s1_readdata),        //                                                                .readdata
		.sys_gpio_bd_s1_writedata                                              (mm_interconnect_0_sys_gpio_bd_s1_writedata),       //                                                                .writedata
		.sys_gpio_bd_s1_chipselect                                             (mm_interconnect_0_sys_gpio_bd_s1_chipselect),      //                                                                .chipselect
		.sys_gpio_in_s1_address                                                (mm_interconnect_0_sys_gpio_in_s1_address),         //                                                  sys_gpio_in_s1.address
		.sys_gpio_in_s1_write                                                  (mm_interconnect_0_sys_gpio_in_s1_write),           //                                                                .write
		.sys_gpio_in_s1_readdata                                               (mm_interconnect_0_sys_gpio_in_s1_readdata),        //                                                                .readdata
		.sys_gpio_in_s1_writedata                                              (mm_interconnect_0_sys_gpio_in_s1_writedata),       //                                                                .writedata
		.sys_gpio_in_s1_chipselect                                             (mm_interconnect_0_sys_gpio_in_s1_chipselect),      //                                                                .chipselect
		.sys_gpio_out_s1_address                                               (mm_interconnect_0_sys_gpio_out_s1_address),        //                                                 sys_gpio_out_s1.address
		.sys_gpio_out_s1_write                                                 (mm_interconnect_0_sys_gpio_out_s1_write),          //                                                                .write
		.sys_gpio_out_s1_readdata                                              (mm_interconnect_0_sys_gpio_out_s1_readdata),       //                                                                .readdata
		.sys_gpio_out_s1_writedata                                             (mm_interconnect_0_sys_gpio_out_s1_writedata),      //                                                                .writedata
		.sys_gpio_out_s1_chipselect                                            (mm_interconnect_0_sys_gpio_out_s1_chipselect),     //                                                                .chipselect
		.sys_id_control_slave_address                                          (mm_interconnect_0_sys_id_control_slave_address),   //                                            sys_id_control_slave.address
		.sys_id_control_slave_readdata                                         (mm_interconnect_0_sys_id_control_slave_readdata)   //                                                                .readdata
	);

	system_bd_mm_interconnect_1 mm_interconnect_1 (
		.spi_dmac_0_m_dest_axi_awid                                         (spi_dmac_0_m_dest_axi_awid),                        //                                        spi_dmac_0_m_dest_axi.awid
		.spi_dmac_0_m_dest_axi_awaddr                                       (spi_dmac_0_m_dest_axi_awaddr),                      //                                                             .awaddr
		.spi_dmac_0_m_dest_axi_awlen                                        (spi_dmac_0_m_dest_axi_awlen),                       //                                                             .awlen
		.spi_dmac_0_m_dest_axi_awsize                                       (spi_dmac_0_m_dest_axi_awsize),                      //                                                             .awsize
		.spi_dmac_0_m_dest_axi_awburst                                      (spi_dmac_0_m_dest_axi_awburst),                     //                                                             .awburst
		.spi_dmac_0_m_dest_axi_awlock                                       (spi_dmac_0_m_dest_axi_awlock),                      //                                                             .awlock
		.spi_dmac_0_m_dest_axi_awcache                                      (spi_dmac_0_m_dest_axi_awcache),                     //                                                             .awcache
		.spi_dmac_0_m_dest_axi_awprot                                       (spi_dmac_0_m_dest_axi_awprot),                      //                                                             .awprot
		.spi_dmac_0_m_dest_axi_awvalid                                      (spi_dmac_0_m_dest_axi_awvalid),                     //                                                             .awvalid
		.spi_dmac_0_m_dest_axi_awready                                      (spi_dmac_0_m_dest_axi_awready),                     //                                                             .awready
		.spi_dmac_0_m_dest_axi_wid                                          (spi_dmac_0_m_dest_axi_wid),                         //                                                             .wid
		.spi_dmac_0_m_dest_axi_wdata                                        (spi_dmac_0_m_dest_axi_wdata),                       //                                                             .wdata
		.spi_dmac_0_m_dest_axi_wstrb                                        (spi_dmac_0_m_dest_axi_wstrb),                       //                                                             .wstrb
		.spi_dmac_0_m_dest_axi_wlast                                        (spi_dmac_0_m_dest_axi_wlast),                       //                                                             .wlast
		.spi_dmac_0_m_dest_axi_wvalid                                       (spi_dmac_0_m_dest_axi_wvalid),                      //                                                             .wvalid
		.spi_dmac_0_m_dest_axi_wready                                       (spi_dmac_0_m_dest_axi_wready),                      //                                                             .wready
		.spi_dmac_0_m_dest_axi_bid                                          (spi_dmac_0_m_dest_axi_bid),                         //                                                             .bid
		.spi_dmac_0_m_dest_axi_bresp                                        (spi_dmac_0_m_dest_axi_bresp),                       //                                                             .bresp
		.spi_dmac_0_m_dest_axi_bvalid                                       (spi_dmac_0_m_dest_axi_bvalid),                      //                                                             .bvalid
		.spi_dmac_0_m_dest_axi_bready                                       (spi_dmac_0_m_dest_axi_bready),                      //                                                             .bready
		.spi_dmac_0_m_dest_axi_arid                                         (spi_dmac_0_m_dest_axi_arid),                        //                                                             .arid
		.spi_dmac_0_m_dest_axi_araddr                                       (spi_dmac_0_m_dest_axi_araddr),                      //                                                             .araddr
		.spi_dmac_0_m_dest_axi_arlen                                        (spi_dmac_0_m_dest_axi_arlen),                       //                                                             .arlen
		.spi_dmac_0_m_dest_axi_arsize                                       (spi_dmac_0_m_dest_axi_arsize),                      //                                                             .arsize
		.spi_dmac_0_m_dest_axi_arburst                                      (spi_dmac_0_m_dest_axi_arburst),                     //                                                             .arburst
		.spi_dmac_0_m_dest_axi_arlock                                       (spi_dmac_0_m_dest_axi_arlock),                      //                                                             .arlock
		.spi_dmac_0_m_dest_axi_arcache                                      (spi_dmac_0_m_dest_axi_arcache),                     //                                                             .arcache
		.spi_dmac_0_m_dest_axi_arprot                                       (spi_dmac_0_m_dest_axi_arprot),                      //                                                             .arprot
		.spi_dmac_0_m_dest_axi_arvalid                                      (spi_dmac_0_m_dest_axi_arvalid),                     //                                                             .arvalid
		.spi_dmac_0_m_dest_axi_arready                                      (spi_dmac_0_m_dest_axi_arready),                     //                                                             .arready
		.spi_dmac_0_m_dest_axi_rid                                          (spi_dmac_0_m_dest_axi_rid),                         //                                                             .rid
		.spi_dmac_0_m_dest_axi_rdata                                        (spi_dmac_0_m_dest_axi_rdata),                       //                                                             .rdata
		.spi_dmac_0_m_dest_axi_rresp                                        (spi_dmac_0_m_dest_axi_rresp),                       //                                                             .rresp
		.spi_dmac_0_m_dest_axi_rlast                                        (spi_dmac_0_m_dest_axi_rlast),                       //                                                             .rlast
		.spi_dmac_0_m_dest_axi_rvalid                                       (spi_dmac_0_m_dest_axi_rvalid),                      //                                                             .rvalid
		.spi_dmac_0_m_dest_axi_rready                                       (spi_dmac_0_m_dest_axi_rready),                      //                                                             .rready
		.sys_hps_f2h_sdram1_data_awid                                       (mm_interconnect_1_sys_hps_f2h_sdram1_data_awid),    //                                      sys_hps_f2h_sdram1_data.awid
		.sys_hps_f2h_sdram1_data_awaddr                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_awaddr),  //                                                             .awaddr
		.sys_hps_f2h_sdram1_data_awlen                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_awlen),   //                                                             .awlen
		.sys_hps_f2h_sdram1_data_awsize                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_awsize),  //                                                             .awsize
		.sys_hps_f2h_sdram1_data_awburst                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_awburst), //                                                             .awburst
		.sys_hps_f2h_sdram1_data_awlock                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_awlock),  //                                                             .awlock
		.sys_hps_f2h_sdram1_data_awcache                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_awcache), //                                                             .awcache
		.sys_hps_f2h_sdram1_data_awprot                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_awprot),  //                                                             .awprot
		.sys_hps_f2h_sdram1_data_awvalid                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_awvalid), //                                                             .awvalid
		.sys_hps_f2h_sdram1_data_awready                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_awready), //                                                             .awready
		.sys_hps_f2h_sdram1_data_wid                                        (mm_interconnect_1_sys_hps_f2h_sdram1_data_wid),     //                                                             .wid
		.sys_hps_f2h_sdram1_data_wdata                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_wdata),   //                                                             .wdata
		.sys_hps_f2h_sdram1_data_wstrb                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_wstrb),   //                                                             .wstrb
		.sys_hps_f2h_sdram1_data_wlast                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_wlast),   //                                                             .wlast
		.sys_hps_f2h_sdram1_data_wvalid                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_wvalid),  //                                                             .wvalid
		.sys_hps_f2h_sdram1_data_wready                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_wready),  //                                                             .wready
		.sys_hps_f2h_sdram1_data_bid                                        (mm_interconnect_1_sys_hps_f2h_sdram1_data_bid),     //                                                             .bid
		.sys_hps_f2h_sdram1_data_bresp                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_bresp),   //                                                             .bresp
		.sys_hps_f2h_sdram1_data_bvalid                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_bvalid),  //                                                             .bvalid
		.sys_hps_f2h_sdram1_data_bready                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_bready),  //                                                             .bready
		.sys_hps_f2h_sdram1_data_arid                                       (mm_interconnect_1_sys_hps_f2h_sdram1_data_arid),    //                                                             .arid
		.sys_hps_f2h_sdram1_data_araddr                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_araddr),  //                                                             .araddr
		.sys_hps_f2h_sdram1_data_arlen                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_arlen),   //                                                             .arlen
		.sys_hps_f2h_sdram1_data_arsize                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_arsize),  //                                                             .arsize
		.sys_hps_f2h_sdram1_data_arburst                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_arburst), //                                                             .arburst
		.sys_hps_f2h_sdram1_data_arlock                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_arlock),  //                                                             .arlock
		.sys_hps_f2h_sdram1_data_arcache                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_arcache), //                                                             .arcache
		.sys_hps_f2h_sdram1_data_arprot                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_arprot),  //                                                             .arprot
		.sys_hps_f2h_sdram1_data_arvalid                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_arvalid), //                                                             .arvalid
		.sys_hps_f2h_sdram1_data_arready                                    (mm_interconnect_1_sys_hps_f2h_sdram1_data_arready), //                                                             .arready
		.sys_hps_f2h_sdram1_data_rid                                        (mm_interconnect_1_sys_hps_f2h_sdram1_data_rid),     //                                                             .rid
		.sys_hps_f2h_sdram1_data_rdata                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_rdata),   //                                                             .rdata
		.sys_hps_f2h_sdram1_data_rresp                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_rresp),   //                                                             .rresp
		.sys_hps_f2h_sdram1_data_rlast                                      (mm_interconnect_1_sys_hps_f2h_sdram1_data_rlast),   //                                                             .rlast
		.sys_hps_f2h_sdram1_data_rvalid                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_rvalid),  //                                                             .rvalid
		.sys_hps_f2h_sdram1_data_rready                                     (mm_interconnect_1_sys_hps_f2h_sdram1_data_rready),  //                                                             .rready
		.sys_hps_h2f_user1_clock_clk                                        (sys_hps_h2f_user1_clock_clk),                       //                                      sys_hps_h2f_user1_clock.clk
		.spi_dmac_0_m_dest_axi_id_pad_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                // spi_dmac_0_m_dest_axi_id_pad_clk_reset_reset_bridge_in_reset.reset
		.spi_dmac_0_m_dest_axi_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset)                     //            spi_dmac_0_m_dest_axi_reset_reset_bridge_in_reset.reset
	);

	system_bd_mm_interconnect_2 mm_interconnect_2 (
		.hdmi_dmac_0_m_src_axi_awid                                           (hdmi_dmac_0_m_src_axi_awid),                              //                                          hdmi_dmac_0_m_src_axi.awid
		.hdmi_dmac_0_m_src_axi_awaddr                                         (hdmi_dmac_0_m_src_axi_awaddr),                            //                                                               .awaddr
		.hdmi_dmac_0_m_src_axi_awlen                                          (hdmi_dmac_0_m_src_axi_awlen),                             //                                                               .awlen
		.hdmi_dmac_0_m_src_axi_awsize                                         (hdmi_dmac_0_m_src_axi_awsize),                            //                                                               .awsize
		.hdmi_dmac_0_m_src_axi_awburst                                        (hdmi_dmac_0_m_src_axi_awburst),                           //                                                               .awburst
		.hdmi_dmac_0_m_src_axi_awlock                                         (hdmi_dmac_0_m_src_axi_awlock),                            //                                                               .awlock
		.hdmi_dmac_0_m_src_axi_awcache                                        (hdmi_dmac_0_m_src_axi_awcache),                           //                                                               .awcache
		.hdmi_dmac_0_m_src_axi_awprot                                         (hdmi_dmac_0_m_src_axi_awprot),                            //                                                               .awprot
		.hdmi_dmac_0_m_src_axi_awvalid                                        (hdmi_dmac_0_m_src_axi_awvalid),                           //                                                               .awvalid
		.hdmi_dmac_0_m_src_axi_awready                                        (hdmi_dmac_0_m_src_axi_awready),                           //                                                               .awready
		.hdmi_dmac_0_m_src_axi_wid                                            (hdmi_dmac_0_m_src_axi_wid),                               //                                                               .wid
		.hdmi_dmac_0_m_src_axi_wdata                                          (hdmi_dmac_0_m_src_axi_wdata),                             //                                                               .wdata
		.hdmi_dmac_0_m_src_axi_wstrb                                          (hdmi_dmac_0_m_src_axi_wstrb),                             //                                                               .wstrb
		.hdmi_dmac_0_m_src_axi_wlast                                          (hdmi_dmac_0_m_src_axi_wlast),                             //                                                               .wlast
		.hdmi_dmac_0_m_src_axi_wvalid                                         (hdmi_dmac_0_m_src_axi_wvalid),                            //                                                               .wvalid
		.hdmi_dmac_0_m_src_axi_wready                                         (hdmi_dmac_0_m_src_axi_wready),                            //                                                               .wready
		.hdmi_dmac_0_m_src_axi_bid                                            (hdmi_dmac_0_m_src_axi_bid),                               //                                                               .bid
		.hdmi_dmac_0_m_src_axi_bresp                                          (hdmi_dmac_0_m_src_axi_bresp),                             //                                                               .bresp
		.hdmi_dmac_0_m_src_axi_bvalid                                         (hdmi_dmac_0_m_src_axi_bvalid),                            //                                                               .bvalid
		.hdmi_dmac_0_m_src_axi_bready                                         (hdmi_dmac_0_m_src_axi_bready),                            //                                                               .bready
		.hdmi_dmac_0_m_src_axi_arid                                           (hdmi_dmac_0_m_src_axi_arid),                              //                                                               .arid
		.hdmi_dmac_0_m_src_axi_araddr                                         (hdmi_dmac_0_m_src_axi_araddr),                            //                                                               .araddr
		.hdmi_dmac_0_m_src_axi_arlen                                          (hdmi_dmac_0_m_src_axi_arlen),                             //                                                               .arlen
		.hdmi_dmac_0_m_src_axi_arsize                                         (hdmi_dmac_0_m_src_axi_arsize),                            //                                                               .arsize
		.hdmi_dmac_0_m_src_axi_arburst                                        (hdmi_dmac_0_m_src_axi_arburst),                           //                                                               .arburst
		.hdmi_dmac_0_m_src_axi_arlock                                         (hdmi_dmac_0_m_src_axi_arlock),                            //                                                               .arlock
		.hdmi_dmac_0_m_src_axi_arcache                                        (hdmi_dmac_0_m_src_axi_arcache),                           //                                                               .arcache
		.hdmi_dmac_0_m_src_axi_arprot                                         (hdmi_dmac_0_m_src_axi_arprot),                            //                                                               .arprot
		.hdmi_dmac_0_m_src_axi_arvalid                                        (hdmi_dmac_0_m_src_axi_arvalid),                           //                                                               .arvalid
		.hdmi_dmac_0_m_src_axi_arready                                        (hdmi_dmac_0_m_src_axi_arready),                           //                                                               .arready
		.hdmi_dmac_0_m_src_axi_rid                                            (hdmi_dmac_0_m_src_axi_rid),                               //                                                               .rid
		.hdmi_dmac_0_m_src_axi_rdata                                          (hdmi_dmac_0_m_src_axi_rdata),                             //                                                               .rdata
		.hdmi_dmac_0_m_src_axi_rresp                                          (hdmi_dmac_0_m_src_axi_rresp),                             //                                                               .rresp
		.hdmi_dmac_0_m_src_axi_rlast                                          (hdmi_dmac_0_m_src_axi_rlast),                             //                                                               .rlast
		.hdmi_dmac_0_m_src_axi_rvalid                                         (hdmi_dmac_0_m_src_axi_rvalid),                            //                                                               .rvalid
		.hdmi_dmac_0_m_src_axi_rready                                         (hdmi_dmac_0_m_src_axi_rready),                            //                                                               .rready
		.sys_hps_h2f_user1_clock_clk                                          (sys_hps_h2f_user1_clock_clk),                             //                                        sys_hps_h2f_user1_clock.clk
		.hdmi_dmac_0_m_src_axi_reset_reset_bridge_in_reset_reset              (rst_controller_reset_out_reset),                          //              hdmi_dmac_0_m_src_axi_reset_reset_bridge_in_reset.reset
		.sys_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                      // sys_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.sys_hps_f2h_sdram0_data_address                                      (mm_interconnect_2_sys_hps_f2h_sdram0_data_address),       //                                        sys_hps_f2h_sdram0_data.address
		.sys_hps_f2h_sdram0_data_write                                        (mm_interconnect_2_sys_hps_f2h_sdram0_data_write),         //                                                               .write
		.sys_hps_f2h_sdram0_data_read                                         (mm_interconnect_2_sys_hps_f2h_sdram0_data_read),          //                                                               .read
		.sys_hps_f2h_sdram0_data_readdata                                     (mm_interconnect_2_sys_hps_f2h_sdram0_data_readdata),      //                                                               .readdata
		.sys_hps_f2h_sdram0_data_writedata                                    (mm_interconnect_2_sys_hps_f2h_sdram0_data_writedata),     //                                                               .writedata
		.sys_hps_f2h_sdram0_data_burstcount                                   (mm_interconnect_2_sys_hps_f2h_sdram0_data_burstcount),    //                                                               .burstcount
		.sys_hps_f2h_sdram0_data_byteenable                                   (mm_interconnect_2_sys_hps_f2h_sdram0_data_byteenable),    //                                                               .byteenable
		.sys_hps_f2h_sdram0_data_readdatavalid                                (mm_interconnect_2_sys_hps_f2h_sdram0_data_readdatavalid), //                                                               .readdatavalid
		.sys_hps_f2h_sdram0_data_waitrequest                                  (mm_interconnect_2_sys_hps_f2h_sdram0_data_waitrequest)    //                                                               .waitrequest
	);

	system_bd_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq), // receiver4.irq
		.sender_irq    (sys_hps_f2h_irq0_irq)      //    sender.irq
	);

	system_bd_irq_mapper_001 irq_mapper_001 (
		.clk        (),                     //       clk.clk
		.reset      (),                     // clk_reset.reset
		.sender_irq (sys_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~sys_rst_reset_n),               // reset_in0.reset
		.clk            (sys_hps_h2f_user1_clock_clk),    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~sys_hps_h2f_reset_reset_n),         // reset_in0.reset
		.clk            (sys_hps_h2f_user1_clock_clk),        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
