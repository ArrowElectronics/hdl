
module clk1 (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
