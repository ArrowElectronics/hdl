// system_bd.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module system_bd (
		inout  wire [19:0] adrv9001_gpio_export,                    //     adrv9001_gpio.export
		input  wire        adrv9001_if_rx1_dclk_in_p_dclk_in,       //       adrv9001_if.rx1_dclk_in_p_dclk_in
		input  wire        adrv9001_if_rx1_idata_in_n_idata0,       //                  .rx1_idata_in_n_idata0
		input  wire        adrv9001_if_rx1_idata_in_p_idata1,       //                  .rx1_idata_in_p_idata1
		input  wire        adrv9001_if_rx1_qdata_in_n_qdata2,       //                  .rx1_qdata_in_n_qdata2
		input  wire        adrv9001_if_rx1_qdata_in_p_qdata3,       //                  .rx1_qdata_in_p_qdata3
		input  wire        adrv9001_if_rx1_strobe_in_p_strobe_in,   //                  .rx1_strobe_in_p_strobe_in
		output wire        adrv9001_if_rx1_enable,                  //                  .rx1_enable
		input  wire        adrv9001_if_rx2_dclk_in_p_dclk_in,       //                  .rx2_dclk_in_p_dclk_in
		input  wire        adrv9001_if_rx2_idata_in_n_idata0,       //                  .rx2_idata_in_n_idata0
		input  wire        adrv9001_if_rx2_idata_in_p_idata1,       //                  .rx2_idata_in_p_idata1
		input  wire        adrv9001_if_rx2_qdata_in_n_qdata2,       //                  .rx2_qdata_in_n_qdata2
		input  wire        adrv9001_if_rx2_qdata_in_p_qdata3,       //                  .rx2_qdata_in_p_qdata3
		input  wire        adrv9001_if_rx2_strobe_in_p_strobe_in,   //                  .rx2_strobe_in_p_strobe_in
		output wire        adrv9001_if_rx2_enable,                  //                  .rx2_enable
		output wire        adrv9001_if_tx1_dclk_out_p_dclk_out,     //                  .tx1_dclk_out_p_dclk_out
		input  wire        adrv9001_if_tx1_dclk_in_p_dclk_in,       //                  .tx1_dclk_in_p_dclk_in
		output wire        adrv9001_if_tx1_idata_out_n_idata0,      //                  .tx1_idata_out_n_idata0
		output wire        adrv9001_if_tx1_idata_out_p_idata1,      //                  .tx1_idata_out_p_idata1
		output wire        adrv9001_if_tx1_qdata_out_n_qdata2,      //                  .tx1_qdata_out_n_qdata2
		output wire        adrv9001_if_tx1_qdata_out_p_qdata3,      //                  .tx1_qdata_out_p_qdata3
		output wire        adrv9001_if_tx1_strobe_out_p_strobe_out, //                  .tx1_strobe_out_p_strobe_out
		output wire        adrv9001_if_tx1_enable,                  //                  .tx1_enable
		output wire        adrv9001_if_tx2_dclk_out_p_dclk_out,     //                  .tx2_dclk_out_p_dclk_out
		input  wire        adrv9001_if_tx2_dclk_in_p_dclk_in,       //                  .tx2_dclk_in_p_dclk_in
		output wire        adrv9001_if_tx2_idata_out_n_idata0,      //                  .tx2_idata_out_n_idata0
		output wire        adrv9001_if_tx2_idata_out_p_idata1,      //                  .tx2_idata_out_p_idata1
		output wire        adrv9001_if_tx2_qdata_out_n_qdata2,      //                  .tx2_qdata_out_n_qdata2
		output wire        adrv9001_if_tx2_qdata_out_p_qdata3,      //                  .tx2_qdata_out_p_qdata3
		output wire        adrv9001_if_tx2_strobe_out_p_strobe_out, //                  .tx2_strobe_out_p_strobe_out
		output wire        adrv9001_if_tx2_enable,                  //                  .tx2_enable
		input  wire        adrv9001_tdd_if_rx1_enable_in,           //   adrv9001_tdd_if.rx1_enable_in
		input  wire        adrv9001_tdd_if_rx2_enable_in,           //                  .rx2_enable_in
		input  wire        adrv9001_tdd_if_tx1_enable_in,           //                  .tx1_enable_in
		input  wire        adrv9001_tdd_if_tx2_enable_in,           //                  .tx2_enable_in
		input  wire        adrv9001_tdd_if_tdd_sync_in,             //                  .tdd_sync_in
		output wire        hdmi_out_h_clk,                          //          hdmi_out.h_clk
		output wire        hdmi_out_h16_hsync,                      //                  .h16_hsync
		output wire        hdmi_out_h16_vsync,                      //                  .h16_vsync
		output wire        hdmi_out_h16_data_e,                     //                  .h16_data_e
		output wire [15:0] hdmi_out_h16_data,                       //                  .h16_data
		output wire [15:0] hdmi_out_h16_es_data,                    //                  .h16_es_data
		output wire        hdmi_out_h24_hsync,                      //                  .h24_hsync
		output wire        hdmi_out_h24_vsync,                      //                  .h24_vsync
		output wire        hdmi_out_h24_data_e,                     //                  .h24_data_e
		output wire [23:0] hdmi_out_h24_data,                       //                  .h24_data
		output wire        hdmi_out_h36_hsync,                      //                  .h36_hsync
		output wire        hdmi_out_h36_vsync,                      //                  .h36_vsync
		output wire        hdmi_out_h36_data_e,                     //                  .h36_data_e
		output wire [35:0] hdmi_out_h36_data,                       //                  .h36_data
		input  wire        spi_0_external_MISO,                     //    spi_0_external.MISO
		output wire        spi_0_external_MOSI,                     //                  .MOSI
		output wire        spi_0_external_SCLK,                     //                  .SCLK
		output wire        spi_0_external_SS_n,                     //                  .SS_n
		input  wire        sys_clk_clk,                             //           sys_clk.clk
		input  wire [31:0] sys_gpio_bd_in_port,                     //       sys_gpio_bd.in_port
		output wire [31:0] sys_gpio_bd_out_port,                    //                  .out_port
		input  wire [31:0] sys_gpio_in_export,                      //       sys_gpio_in.export
		output wire [31:0] sys_gpio_out_export,                     //      sys_gpio_out.export
		output wire        sys_hps_h2f_reset_reset_n,               // sys_hps_h2f_reset.reset_n
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TX_CLK, //    sys_hps_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD0,   //                  .hps_io_emac1_inst_TXD0
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD1,   //                  .hps_io_emac1_inst_TXD1
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD2,   //                  .hps_io_emac1_inst_TXD2
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TXD3,   //                  .hps_io_emac1_inst_TXD3
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD0,   //                  .hps_io_emac1_inst_RXD0
		inout  wire        sys_hps_hps_io_hps_io_emac1_inst_MDIO,   //                  .hps_io_emac1_inst_MDIO
		output wire        sys_hps_hps_io_hps_io_emac1_inst_MDC,    //                  .hps_io_emac1_inst_MDC
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RX_CTL, //                  .hps_io_emac1_inst_RX_CTL
		output wire        sys_hps_hps_io_hps_io_emac1_inst_TX_CTL, //                  .hps_io_emac1_inst_TX_CTL
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RX_CLK, //                  .hps_io_emac1_inst_RX_CLK
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD1,   //                  .hps_io_emac1_inst_RXD1
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD2,   //                  .hps_io_emac1_inst_RXD2
		input  wire        sys_hps_hps_io_hps_io_emac1_inst_RXD3,   //                  .hps_io_emac1_inst_RXD3
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO0,     //                  .hps_io_qspi_inst_IO0
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO1,     //                  .hps_io_qspi_inst_IO1
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO2,     //                  .hps_io_qspi_inst_IO2
		inout  wire        sys_hps_hps_io_hps_io_qspi_inst_IO3,     //                  .hps_io_qspi_inst_IO3
		output wire        sys_hps_hps_io_hps_io_qspi_inst_SS0,     //                  .hps_io_qspi_inst_SS0
		output wire        sys_hps_hps_io_hps_io_qspi_inst_CLK,     //                  .hps_io_qspi_inst_CLK
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_CMD,     //                  .hps_io_sdio_inst_CMD
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D0,      //                  .hps_io_sdio_inst_D0
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D1,      //                  .hps_io_sdio_inst_D1
		output wire        sys_hps_hps_io_hps_io_sdio_inst_CLK,     //                  .hps_io_sdio_inst_CLK
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D2,      //                  .hps_io_sdio_inst_D2
		inout  wire        sys_hps_hps_io_hps_io_sdio_inst_D3,      //                  .hps_io_sdio_inst_D3
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D0,      //                  .hps_io_usb1_inst_D0
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D1,      //                  .hps_io_usb1_inst_D1
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D2,      //                  .hps_io_usb1_inst_D2
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D3,      //                  .hps_io_usb1_inst_D3
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D4,      //                  .hps_io_usb1_inst_D4
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D5,      //                  .hps_io_usb1_inst_D5
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D6,      //                  .hps_io_usb1_inst_D6
		inout  wire        sys_hps_hps_io_hps_io_usb1_inst_D7,      //                  .hps_io_usb1_inst_D7
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_CLK,     //                  .hps_io_usb1_inst_CLK
		output wire        sys_hps_hps_io_hps_io_usb1_inst_STP,     //                  .hps_io_usb1_inst_STP
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_DIR,     //                  .hps_io_usb1_inst_DIR
		input  wire        sys_hps_hps_io_hps_io_usb1_inst_NXT,     //                  .hps_io_usb1_inst_NXT
		input  wire        sys_hps_hps_io_hps_io_uart0_inst_RX,     //                  .hps_io_uart0_inst_RX
		output wire        sys_hps_hps_io_hps_io_uart0_inst_TX,     //                  .hps_io_uart0_inst_TX
		inout  wire        sys_hps_hps_io_hps_io_i2c0_inst_SDA,     //                  .hps_io_i2c0_inst_SDA
		inout  wire        sys_hps_hps_io_hps_io_i2c0_inst_SCL,     //                  .hps_io_i2c0_inst_SCL
		inout  wire        sys_hps_hps_io_hps_io_i2c1_inst_SDA,     //                  .hps_io_i2c1_inst_SDA
		inout  wire        sys_hps_hps_io_hps_io_i2c1_inst_SCL,     //                  .hps_io_i2c1_inst_SCL
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO00,  //                  .hps_io_gpio_inst_GPIO00
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO09,  //                  .hps_io_gpio_inst_GPIO09
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO35,  //                  .hps_io_gpio_inst_GPIO35
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO40,  //                  .hps_io_gpio_inst_GPIO40
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO41,  //                  .hps_io_gpio_inst_GPIO41
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO42,  //                  .hps_io_gpio_inst_GPIO42
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO43,  //                  .hps_io_gpio_inst_GPIO43
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO44,  //                  .hps_io_gpio_inst_GPIO44
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO48,  //                  .hps_io_gpio_inst_GPIO48
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO53,  //                  .hps_io_gpio_inst_GPIO53
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO54,  //                  .hps_io_gpio_inst_GPIO54
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO55,  //                  .hps_io_gpio_inst_GPIO55
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO56,  //                  .hps_io_gpio_inst_GPIO56
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO57,  //                  .hps_io_gpio_inst_GPIO57
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO58,  //                  .hps_io_gpio_inst_GPIO58
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO59,  //                  .hps_io_gpio_inst_GPIO59
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO61,  //                  .hps_io_gpio_inst_GPIO61
		inout  wire        sys_hps_hps_io_hps_io_gpio_inst_GPIO65,  //                  .hps_io_gpio_inst_GPIO65
		output wire [14:0] sys_hps_memory_mem_a,                    //    sys_hps_memory.mem_a
		output wire [2:0]  sys_hps_memory_mem_ba,                   //                  .mem_ba
		output wire        sys_hps_memory_mem_ck,                   //                  .mem_ck
		output wire        sys_hps_memory_mem_ck_n,                 //                  .mem_ck_n
		output wire        sys_hps_memory_mem_cke,                  //                  .mem_cke
		output wire        sys_hps_memory_mem_cs_n,                 //                  .mem_cs_n
		output wire        sys_hps_memory_mem_ras_n,                //                  .mem_ras_n
		output wire        sys_hps_memory_mem_cas_n,                //                  .mem_cas_n
		output wire        sys_hps_memory_mem_we_n,                 //                  .mem_we_n
		output wire        sys_hps_memory_mem_reset_n,              //                  .mem_reset_n
		inout  wire [31:0] sys_hps_memory_mem_dq,                   //                  .mem_dq
		inout  wire [3:0]  sys_hps_memory_mem_dqs,                  //                  .mem_dqs
		inout  wire [3:0]  sys_hps_memory_mem_dqs_n,                //                  .mem_dqs_n
		output wire        sys_hps_memory_mem_odt,                  //                  .mem_odt
		output wire [3:0]  sys_hps_memory_mem_dm,                   //                  .mem_dm
		input  wire        sys_hps_memory_oct_rzqin,                //                  .oct_rzqin
		input  wire        sys_rst_reset_n                          //           sys_rst.reset_n
	);

	wire         axi_dac_dma_m_axis_tvalid;                               // axi_dac_dma:m_axis_valid -> util_dac_upack:s_axis_valid
	wire         axi_dac_dma_m_axis_tready;                               // util_dac_upack:s_axis_ready -> axi_dac_dma:m_axis_ready
	wire  [63:0] axi_dac_dma_m_axis_tdata;                                // axi_dac_dma:m_axis_data -> util_dac_upack:s_axis_data
	wire         hdmi_dmac_0_m_axis_tvalid;                               // hdmi_dmac_0:m_axis_valid -> axi_hdmi_tx_0:vdma_valid
	wire         hdmi_dmac_0_m_axis_tready;                               // axi_hdmi_tx_0:vdma_ready -> hdmi_dmac_0:m_axis_ready
	wire         hdmi_dmac_0_m_axis_tlast;                                // hdmi_dmac_0:m_axis_last -> axi_hdmi_tx_0:vdma_end_of_frame
	wire  [63:0] hdmi_dmac_0_m_axis_tdata;                                // hdmi_dmac_0:m_axis_data -> axi_hdmi_tx_0:vdma_data
	wire         sys_hps_h2f_user1_clock_clk;                             // sys_hps:h2f_user1_clk -> [avl_adrv9001_gpio:clk, axi_adc_dma:fifo_wr_clk, axi_adc_dma:m_dest_axi_aclk, axi_adc_dma:s_axi_aclk, axi_adrv9001:s_axi_aclk, axi_dac_dma:m_axis_aclk, axi_dac_dma:m_src_axi_aclk, axi_dac_dma:s_axi_aclk, axi_hdmi_tx_0:s_axi_aclk, axi_hdmi_tx_0:vdma_clk, hdmi_dmac_0:m_axis_aclk, hdmi_dmac_0:m_src_axi_aclk, hdmi_dmac_0:s_axi_aclk, hdmi_pll:refclk, mm_interconnect_0:sys_hps_h2f_user1_clock_clk, mm_interconnect_1:sys_hps_h2f_user1_clock_clk, rst_controller:clk, rst_controller_001:clk, spi_0:clk, sys_gpio_bd:clk, sys_gpio_in:clk, sys_gpio_out:clk, sys_hps:f2h_axi_clk, sys_hps:f2h_sdram0_clk, sys_hps:f2h_sdram1_clk, sys_hps:f2h_sdram2_clk, sys_hps:h2f_axi_clk, sys_hps:h2f_lw_axi_clk, sys_id:clock, util_adc_pack:clk, util_adc_wfifo:dout_clk, util_dac_rfifo:din_clk, util_dac_upack:clk]
	wire         axi_adrv9001_if_adc_1_clk_clk;                           // axi_adrv9001:adc_1_clk -> util_adc_wfifo:din_clk
	wire         axi_adrv9001_if_dac_1_clk_clk;                           // axi_adrv9001:dac_1_clk -> util_dac_rfifo:dout_clk
	wire         hdmi_pll_outclk0_clk;                                    // hdmi_pll:outclk_0 -> axi_hdmi_tx_0:hdmi_clk
	wire         axi_adrv9001_adc_1_ch_0_valid;                           // axi_adrv9001:adc_1_valid_i0 -> util_adc_wfifo:din_valid_0
	wire  [15:0] axi_adrv9001_adc_1_ch_0_data;                            // axi_adrv9001:adc_1_data_i0 -> util_adc_wfifo:din_data_0
	wire         axi_adrv9001_adc_1_ch_0_enable;                          // axi_adrv9001:adc_1_enable_i0 -> util_adc_wfifo:din_enable_0
	wire         axi_adrv9001_adc_1_ch_1_valid;                           // axi_adrv9001:adc_1_valid_q0 -> util_adc_wfifo:din_valid_1
	wire  [15:0] axi_adrv9001_adc_1_ch_1_data;                            // axi_adrv9001:adc_1_data_q0 -> util_adc_wfifo:din_data_1
	wire         axi_adrv9001_adc_1_ch_1_enable;                          // axi_adrv9001:adc_1_enable_q0 -> util_adc_wfifo:din_enable_1
	wire         axi_adrv9001_adc_1_ch_2_valid;                           // axi_adrv9001:adc_1_valid_i1 -> util_adc_wfifo:din_valid_2
	wire  [15:0] axi_adrv9001_adc_1_ch_2_data;                            // axi_adrv9001:adc_1_data_i1 -> util_adc_wfifo:din_data_2
	wire         axi_adrv9001_adc_1_ch_2_enable;                          // axi_adrv9001:adc_1_enable_i1 -> util_adc_wfifo:din_enable_2
	wire         axi_adrv9001_adc_1_ch_3_valid;                           // axi_adrv9001:adc_1_valid_q1 -> util_adc_wfifo:din_valid_3
	wire  [15:0] axi_adrv9001_adc_1_ch_3_data;                            // axi_adrv9001:adc_1_data_q1 -> util_adc_wfifo:din_data_3
	wire         axi_adrv9001_adc_1_ch_3_enable;                          // axi_adrv9001:adc_1_enable_q1 -> util_adc_wfifo:din_enable_3
	wire         util_dac_rfifo_din_0_valid;                              // util_dac_rfifo:din_valid_0 -> util_dac_upack:fifo_rd_en_0
	wire  [15:0] util_dac_upack_dac_ch_0_data;                            // util_dac_upack:fifo_rd_data_0 -> util_dac_rfifo:din_data_0
	wire         util_dac_rfifo_din_0_enable;                             // util_dac_rfifo:din_enable_0 -> util_dac_upack:enable_0
	wire         util_dac_upack_dac_ch_0_data_valid;                      // util_dac_upack:fifo_rd_valid_0 -> util_dac_rfifo:din_valid_in_0
	wire         util_dac_rfifo_din_1_valid;                              // util_dac_rfifo:din_valid_1 -> util_dac_upack:fifo_rd_en_1
	wire  [15:0] util_dac_upack_dac_ch_1_data;                            // util_dac_upack:fifo_rd_data_1 -> util_dac_rfifo:din_data_1
	wire         util_dac_rfifo_din_1_enable;                             // util_dac_rfifo:din_enable_1 -> util_dac_upack:enable_1
	wire         util_dac_upack_dac_ch_1_data_valid;                      // util_dac_upack:fifo_rd_valid_1 -> util_dac_rfifo:din_valid_in_1
	wire         util_dac_rfifo_din_2_valid;                              // util_dac_rfifo:din_valid_2 -> util_dac_upack:fifo_rd_en_2
	wire  [15:0] util_dac_upack_dac_ch_2_data;                            // util_dac_upack:fifo_rd_data_2 -> util_dac_rfifo:din_data_2
	wire         util_dac_rfifo_din_2_enable;                             // util_dac_rfifo:din_enable_2 -> util_dac_upack:enable_2
	wire         util_dac_upack_dac_ch_2_data_valid;                      // util_dac_upack:fifo_rd_valid_2 -> util_dac_rfifo:din_valid_in_2
	wire         util_dac_rfifo_din_3_valid;                              // util_dac_rfifo:din_valid_3 -> util_dac_upack:fifo_rd_en_3
	wire  [15:0] util_dac_upack_dac_ch_3_data;                            // util_dac_upack:fifo_rd_data_3 -> util_dac_rfifo:din_data_3
	wire         util_dac_rfifo_din_3_enable;                             // util_dac_rfifo:din_enable_3 -> util_dac_upack:enable_3
	wire         util_dac_upack_dac_ch_3_data_valid;                      // util_dac_upack:fifo_rd_valid_3 -> util_dac_rfifo:din_valid_in_3
	wire         util_adc_wfifo_dout_0_valid;                             // util_adc_wfifo:dout_valid_0 -> util_adc_pack:fifo_wr_en_0
	wire  [15:0] util_adc_wfifo_dout_0_data;                              // util_adc_wfifo:dout_data_0 -> util_adc_pack:fifo_wr_data_0
	wire         util_adc_wfifo_dout_0_enable;                            // util_adc_wfifo:dout_enable_0 -> util_adc_pack:enable_0
	wire         axi_adrv9001_dac_1_ch_0_valid;                           // axi_adrv9001:dac_1_valid_i0 -> util_dac_rfifo:dout_valid_0
	wire  [15:0] util_dac_rfifo_dout_0_data;                              // util_dac_rfifo:dout_data_0 -> axi_adrv9001:dac_1_data_i0
	wire         axi_adrv9001_dac_1_ch_0_enable;                          // axi_adrv9001:dac_1_enable_i0 -> util_dac_rfifo:dout_enable_0
	wire         util_adc_wfifo_dout_1_valid;                             // util_adc_wfifo:dout_valid_1 -> util_adc_pack:fifo_wr_en_1
	wire  [15:0] util_adc_wfifo_dout_1_data;                              // util_adc_wfifo:dout_data_1 -> util_adc_pack:fifo_wr_data_1
	wire         util_adc_wfifo_dout_1_enable;                            // util_adc_wfifo:dout_enable_1 -> util_adc_pack:enable_1
	wire         axi_adrv9001_dac_1_ch_1_valid;                           // axi_adrv9001:dac_1_valid_q0 -> util_dac_rfifo:dout_valid_1
	wire  [15:0] util_dac_rfifo_dout_1_data;                              // util_dac_rfifo:dout_data_1 -> axi_adrv9001:dac_1_data_q0
	wire         axi_adrv9001_dac_1_ch_1_enable;                          // axi_adrv9001:dac_1_enable_q0 -> util_dac_rfifo:dout_enable_1
	wire         util_adc_wfifo_dout_2_valid;                             // util_adc_wfifo:dout_valid_2 -> util_adc_pack:fifo_wr_en_2
	wire  [15:0] util_adc_wfifo_dout_2_data;                              // util_adc_wfifo:dout_data_2 -> util_adc_pack:fifo_wr_data_2
	wire         util_adc_wfifo_dout_2_enable;                            // util_adc_wfifo:dout_enable_2 -> util_adc_pack:enable_2
	wire         axi_adrv9001_dac_1_ch_2_valid;                           // axi_adrv9001:dac_1_valid_i1 -> util_dac_rfifo:dout_valid_2
	wire  [15:0] util_dac_rfifo_dout_2_data;                              // util_dac_rfifo:dout_data_2 -> axi_adrv9001:dac_1_data_i1
	wire         axi_adrv9001_dac_1_ch_2_enable;                          // axi_adrv9001:dac_1_enable_i1 -> util_dac_rfifo:dout_enable_2
	wire         util_adc_wfifo_dout_3_valid;                             // util_adc_wfifo:dout_valid_3 -> util_adc_pack:fifo_wr_en_3
	wire  [15:0] util_adc_wfifo_dout_3_data;                              // util_adc_wfifo:dout_data_3 -> util_adc_pack:fifo_wr_data_3
	wire         util_adc_wfifo_dout_3_enable;                            // util_adc_wfifo:dout_enable_3 -> util_adc_pack:enable_3
	wire         axi_adrv9001_dac_1_ch_3_valid;                           // axi_adrv9001:dac_1_valid_q1 -> util_dac_rfifo:dout_valid_3
	wire  [15:0] util_dac_rfifo_dout_3_data;                              // util_dac_rfifo:dout_data_3 -> axi_adrv9001:dac_1_data_q1
	wire         axi_adrv9001_dac_1_ch_3_enable;                          // axi_adrv9001:dac_1_enable_q1 -> util_dac_rfifo:dout_enable_3
	wire         util_adc_wfifo_if_din_ovf_ovf;                           // util_adc_wfifo:din_ovf -> axi_adrv9001:adc_1_dovf
	wire         util_dac_rfifo_if_dout_unf_unf;                          // util_dac_rfifo:dout_unf -> axi_adrv9001:dac_1_dunf
	wire         util_dac_upack_if_fifo_rd_underflow_unf;                 // util_dac_upack:fifo_rd_underflow -> util_dac_rfifo:din_unf
	wire         util_adc_pack_if_fifo_wr_overflow_ovf;                   // util_adc_pack:fifo_wr_overflow -> util_adc_wfifo:dout_ovf
	wire         axi_adc_dma_if_fifo_wr_overflow_ovf;                     // axi_adc_dma:fifo_wr_overflow -> util_adc_pack:packed_fifo_wr_overflow
	wire  [63:0] util_adc_pack_if_packed_fifo_wr_data_data;               // util_adc_pack:packed_fifo_wr_data -> axi_adc_dma:fifo_wr_din
	wire         util_adc_pack_if_packed_fifo_wr_en_valid;                // util_adc_pack:packed_fifo_wr_en -> axi_adc_dma:fifo_wr_en
	wire         util_adc_pack_if_packed_fifo_wr_sync_sync;               // util_adc_pack:packed_fifo_wr_sync -> axi_adc_dma:fifo_wr_sync
	wire         axi_adrv9001_if_adc_1_rst_reset;                         // axi_adrv9001:adc_1_rst -> util_adc_wfifo:din_rst
	wire         axi_adrv9001_if_dac_1_rst_reset;                         // axi_adrv9001:dac_1_rst -> util_dac_rfifo:dout_rst
	wire   [1:0] sys_hps_h2f_lw_axi_master_awburst;                       // sys_hps:h2f_lw_AWBURST -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awburst
	wire   [3:0] sys_hps_h2f_lw_axi_master_arlen;                         // sys_hps:h2f_lw_ARLEN -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arlen
	wire   [3:0] sys_hps_h2f_lw_axi_master_wstrb;                         // sys_hps:h2f_lw_WSTRB -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wstrb
	wire         sys_hps_h2f_lw_axi_master_wready;                        // mm_interconnect_0:sys_hps_h2f_lw_axi_master_wready -> sys_hps:h2f_lw_WREADY
	wire  [11:0] sys_hps_h2f_lw_axi_master_rid;                           // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rid -> sys_hps:h2f_lw_RID
	wire         sys_hps_h2f_lw_axi_master_rready;                        // sys_hps:h2f_lw_RREADY -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_rready
	wire   [3:0] sys_hps_h2f_lw_axi_master_awlen;                         // sys_hps:h2f_lw_AWLEN -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awlen
	wire  [11:0] sys_hps_h2f_lw_axi_master_wid;                           // sys_hps:h2f_lw_WID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wid
	wire   [3:0] sys_hps_h2f_lw_axi_master_arcache;                       // sys_hps:h2f_lw_ARCACHE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arcache
	wire         sys_hps_h2f_lw_axi_master_wvalid;                        // sys_hps:h2f_lw_WVALID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wvalid
	wire  [20:0] sys_hps_h2f_lw_axi_master_araddr;                        // sys_hps:h2f_lw_ARADDR -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_araddr
	wire   [2:0] sys_hps_h2f_lw_axi_master_arprot;                        // sys_hps:h2f_lw_ARPROT -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arprot
	wire   [2:0] sys_hps_h2f_lw_axi_master_awprot;                        // sys_hps:h2f_lw_AWPROT -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awprot
	wire  [31:0] sys_hps_h2f_lw_axi_master_wdata;                         // sys_hps:h2f_lw_WDATA -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wdata
	wire         sys_hps_h2f_lw_axi_master_arvalid;                       // sys_hps:h2f_lw_ARVALID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arvalid
	wire   [3:0] sys_hps_h2f_lw_axi_master_awcache;                       // sys_hps:h2f_lw_AWCACHE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awcache
	wire  [11:0] sys_hps_h2f_lw_axi_master_arid;                          // sys_hps:h2f_lw_ARID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arid
	wire   [1:0] sys_hps_h2f_lw_axi_master_arlock;                        // sys_hps:h2f_lw_ARLOCK -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arlock
	wire   [1:0] sys_hps_h2f_lw_axi_master_awlock;                        // sys_hps:h2f_lw_AWLOCK -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awlock
	wire  [20:0] sys_hps_h2f_lw_axi_master_awaddr;                        // sys_hps:h2f_lw_AWADDR -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awaddr
	wire   [1:0] sys_hps_h2f_lw_axi_master_bresp;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_bresp -> sys_hps:h2f_lw_BRESP
	wire         sys_hps_h2f_lw_axi_master_arready;                       // mm_interconnect_0:sys_hps_h2f_lw_axi_master_arready -> sys_hps:h2f_lw_ARREADY
	wire  [31:0] sys_hps_h2f_lw_axi_master_rdata;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rdata -> sys_hps:h2f_lw_RDATA
	wire         sys_hps_h2f_lw_axi_master_awready;                       // mm_interconnect_0:sys_hps_h2f_lw_axi_master_awready -> sys_hps:h2f_lw_AWREADY
	wire   [1:0] sys_hps_h2f_lw_axi_master_arburst;                       // sys_hps:h2f_lw_ARBURST -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arburst
	wire   [2:0] sys_hps_h2f_lw_axi_master_arsize;                        // sys_hps:h2f_lw_ARSIZE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_arsize
	wire         sys_hps_h2f_lw_axi_master_bready;                        // sys_hps:h2f_lw_BREADY -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_bready
	wire         sys_hps_h2f_lw_axi_master_rlast;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rlast -> sys_hps:h2f_lw_RLAST
	wire         sys_hps_h2f_lw_axi_master_wlast;                         // sys_hps:h2f_lw_WLAST -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_wlast
	wire   [1:0] sys_hps_h2f_lw_axi_master_rresp;                         // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rresp -> sys_hps:h2f_lw_RRESP
	wire  [11:0] sys_hps_h2f_lw_axi_master_awid;                          // sys_hps:h2f_lw_AWID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awid
	wire  [11:0] sys_hps_h2f_lw_axi_master_bid;                           // mm_interconnect_0:sys_hps_h2f_lw_axi_master_bid -> sys_hps:h2f_lw_BID
	wire         sys_hps_h2f_lw_axi_master_bvalid;                        // mm_interconnect_0:sys_hps_h2f_lw_axi_master_bvalid -> sys_hps:h2f_lw_BVALID
	wire   [2:0] sys_hps_h2f_lw_axi_master_awsize;                        // sys_hps:h2f_lw_AWSIZE -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awsize
	wire         sys_hps_h2f_lw_axi_master_awvalid;                       // sys_hps:h2f_lw_AWVALID -> mm_interconnect_0:sys_hps_h2f_lw_axi_master_awvalid
	wire         sys_hps_h2f_lw_axi_master_rvalid;                        // mm_interconnect_0:sys_hps_h2f_lw_axi_master_rvalid -> sys_hps:h2f_lw_RVALID
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;         // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;          // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire         mm_interconnect_0_sys_gpio_bd_s1_chipselect;             // mm_interconnect_0:sys_gpio_bd_s1_chipselect -> sys_gpio_bd:chipselect
	wire  [31:0] mm_interconnect_0_sys_gpio_bd_s1_readdata;               // sys_gpio_bd:readdata -> mm_interconnect_0:sys_gpio_bd_s1_readdata
	wire   [1:0] mm_interconnect_0_sys_gpio_bd_s1_address;                // mm_interconnect_0:sys_gpio_bd_s1_address -> sys_gpio_bd:address
	wire         mm_interconnect_0_sys_gpio_bd_s1_write;                  // mm_interconnect_0:sys_gpio_bd_s1_write -> sys_gpio_bd:write_n
	wire  [31:0] mm_interconnect_0_sys_gpio_bd_s1_writedata;              // mm_interconnect_0:sys_gpio_bd_s1_writedata -> sys_gpio_bd:writedata
	wire         mm_interconnect_0_sys_gpio_in_s1_chipselect;             // mm_interconnect_0:sys_gpio_in_s1_chipselect -> sys_gpio_in:chipselect
	wire  [31:0] mm_interconnect_0_sys_gpio_in_s1_readdata;               // sys_gpio_in:readdata -> mm_interconnect_0:sys_gpio_in_s1_readdata
	wire   [1:0] mm_interconnect_0_sys_gpio_in_s1_address;                // mm_interconnect_0:sys_gpio_in_s1_address -> sys_gpio_in:address
	wire         mm_interconnect_0_sys_gpio_in_s1_write;                  // mm_interconnect_0:sys_gpio_in_s1_write -> sys_gpio_in:write_n
	wire  [31:0] mm_interconnect_0_sys_gpio_in_s1_writedata;              // mm_interconnect_0:sys_gpio_in_s1_writedata -> sys_gpio_in:writedata
	wire         mm_interconnect_0_sys_gpio_out_s1_chipselect;            // mm_interconnect_0:sys_gpio_out_s1_chipselect -> sys_gpio_out:chipselect
	wire  [31:0] mm_interconnect_0_sys_gpio_out_s1_readdata;              // sys_gpio_out:readdata -> mm_interconnect_0:sys_gpio_out_s1_readdata
	wire   [1:0] mm_interconnect_0_sys_gpio_out_s1_address;               // mm_interconnect_0:sys_gpio_out_s1_address -> sys_gpio_out:address
	wire         mm_interconnect_0_sys_gpio_out_s1_write;                 // mm_interconnect_0:sys_gpio_out_s1_write -> sys_gpio_out:write_n
	wire  [31:0] mm_interconnect_0_sys_gpio_out_s1_writedata;             // mm_interconnect_0:sys_gpio_out_s1_writedata -> sys_gpio_out:writedata
	wire         mm_interconnect_0_avl_adrv9001_gpio_s1_chipselect;       // mm_interconnect_0:avl_adrv9001_gpio_s1_chipselect -> avl_adrv9001_gpio:chipselect
	wire  [31:0] mm_interconnect_0_avl_adrv9001_gpio_s1_readdata;         // avl_adrv9001_gpio:readdata -> mm_interconnect_0:avl_adrv9001_gpio_s1_readdata
	wire   [1:0] mm_interconnect_0_avl_adrv9001_gpio_s1_address;          // mm_interconnect_0:avl_adrv9001_gpio_s1_address -> avl_adrv9001_gpio:address
	wire         mm_interconnect_0_avl_adrv9001_gpio_s1_write;            // mm_interconnect_0:avl_adrv9001_gpio_s1_write -> avl_adrv9001_gpio:write_n
	wire  [31:0] mm_interconnect_0_avl_adrv9001_gpio_s1_writedata;        // mm_interconnect_0:avl_adrv9001_gpio_s1_writedata -> avl_adrv9001_gpio:writedata
	wire  [10:0] mm_interconnect_0_hdmi_dmac_0_s_axi_awaddr;              // mm_interconnect_0:hdmi_dmac_0_s_axi_awaddr -> hdmi_dmac_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_hdmi_dmac_0_s_axi_bresp;               // hdmi_dmac_0:s_axi_bresp -> mm_interconnect_0:hdmi_dmac_0_s_axi_bresp
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_arready;             // hdmi_dmac_0:s_axi_arready -> mm_interconnect_0:hdmi_dmac_0_s_axi_arready
	wire  [31:0] mm_interconnect_0_hdmi_dmac_0_s_axi_rdata;               // hdmi_dmac_0:s_axi_rdata -> mm_interconnect_0:hdmi_dmac_0_s_axi_rdata
	wire   [3:0] mm_interconnect_0_hdmi_dmac_0_s_axi_wstrb;               // mm_interconnect_0:hdmi_dmac_0_s_axi_wstrb -> hdmi_dmac_0:s_axi_wstrb
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_wready;              // hdmi_dmac_0:s_axi_wready -> mm_interconnect_0:hdmi_dmac_0_s_axi_wready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_awready;             // hdmi_dmac_0:s_axi_awready -> mm_interconnect_0:hdmi_dmac_0_s_axi_awready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_rready;              // mm_interconnect_0:hdmi_dmac_0_s_axi_rready -> hdmi_dmac_0:s_axi_rready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_bready;              // mm_interconnect_0:hdmi_dmac_0_s_axi_bready -> hdmi_dmac_0:s_axi_bready
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_wvalid;              // mm_interconnect_0:hdmi_dmac_0_s_axi_wvalid -> hdmi_dmac_0:s_axi_wvalid
	wire  [10:0] mm_interconnect_0_hdmi_dmac_0_s_axi_araddr;              // mm_interconnect_0:hdmi_dmac_0_s_axi_araddr -> hdmi_dmac_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_hdmi_dmac_0_s_axi_arprot;              // mm_interconnect_0:hdmi_dmac_0_s_axi_arprot -> hdmi_dmac_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_hdmi_dmac_0_s_axi_rresp;               // hdmi_dmac_0:s_axi_rresp -> mm_interconnect_0:hdmi_dmac_0_s_axi_rresp
	wire   [2:0] mm_interconnect_0_hdmi_dmac_0_s_axi_awprot;              // mm_interconnect_0:hdmi_dmac_0_s_axi_awprot -> hdmi_dmac_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_hdmi_dmac_0_s_axi_wdata;               // mm_interconnect_0:hdmi_dmac_0_s_axi_wdata -> hdmi_dmac_0:s_axi_wdata
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_arvalid;             // mm_interconnect_0:hdmi_dmac_0_s_axi_arvalid -> hdmi_dmac_0:s_axi_arvalid
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_bvalid;              // hdmi_dmac_0:s_axi_bvalid -> mm_interconnect_0:hdmi_dmac_0_s_axi_bvalid
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_awvalid;             // mm_interconnect_0:hdmi_dmac_0_s_axi_awvalid -> hdmi_dmac_0:s_axi_awvalid
	wire         mm_interconnect_0_hdmi_dmac_0_s_axi_rvalid;              // hdmi_dmac_0:s_axi_rvalid -> mm_interconnect_0:hdmi_dmac_0_s_axi_rvalid
	wire  [15:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_awaddr;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_awaddr -> axi_hdmi_tx_0:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_bresp;             // axi_hdmi_tx_0:s_axi_bresp -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_bresp
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_arready;           // axi_hdmi_tx_0:s_axi_arready -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_arready
	wire  [31:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_rdata;             // axi_hdmi_tx_0:s_axi_rdata -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_rdata
	wire   [3:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_wstrb;             // mm_interconnect_0:axi_hdmi_tx_0_s_axi_wstrb -> axi_hdmi_tx_0:s_axi_wstrb
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_wready;            // axi_hdmi_tx_0:s_axi_wready -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_wready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_awready;           // axi_hdmi_tx_0:s_axi_awready -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_awready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_rready;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_rready -> axi_hdmi_tx_0:s_axi_rready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_bready;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_bready -> axi_hdmi_tx_0:s_axi_bready
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_wvalid;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_wvalid -> axi_hdmi_tx_0:s_axi_wvalid
	wire  [15:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_araddr;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_araddr -> axi_hdmi_tx_0:s_axi_araddr
	wire   [2:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_arprot;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_arprot -> axi_hdmi_tx_0:s_axi_arprot
	wire   [1:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_rresp;             // axi_hdmi_tx_0:s_axi_rresp -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_rresp
	wire   [2:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_awprot;            // mm_interconnect_0:axi_hdmi_tx_0_s_axi_awprot -> axi_hdmi_tx_0:s_axi_awprot
	wire  [31:0] mm_interconnect_0_axi_hdmi_tx_0_s_axi_wdata;             // mm_interconnect_0:axi_hdmi_tx_0_s_axi_wdata -> axi_hdmi_tx_0:s_axi_wdata
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_arvalid;           // mm_interconnect_0:axi_hdmi_tx_0_s_axi_arvalid -> axi_hdmi_tx_0:s_axi_arvalid
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_bvalid;            // axi_hdmi_tx_0:s_axi_bvalid -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_bvalid
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_awvalid;           // mm_interconnect_0:axi_hdmi_tx_0_s_axi_awvalid -> axi_hdmi_tx_0:s_axi_awvalid
	wire         mm_interconnect_0_axi_hdmi_tx_0_s_axi_rvalid;            // axi_hdmi_tx_0:s_axi_rvalid -> mm_interconnect_0:axi_hdmi_tx_0_s_axi_rvalid
	wire  [15:0] mm_interconnect_0_axi_adrv9001_s_axi_awaddr;             // mm_interconnect_0:axi_adrv9001_s_axi_awaddr -> axi_adrv9001:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_axi_adrv9001_s_axi_bresp;              // axi_adrv9001:s_axi_bresp -> mm_interconnect_0:axi_adrv9001_s_axi_bresp
	wire         mm_interconnect_0_axi_adrv9001_s_axi_arready;            // axi_adrv9001:s_axi_arready -> mm_interconnect_0:axi_adrv9001_s_axi_arready
	wire  [31:0] mm_interconnect_0_axi_adrv9001_s_axi_rdata;              // axi_adrv9001:s_axi_rdata -> mm_interconnect_0:axi_adrv9001_s_axi_rdata
	wire   [3:0] mm_interconnect_0_axi_adrv9001_s_axi_wstrb;              // mm_interconnect_0:axi_adrv9001_s_axi_wstrb -> axi_adrv9001:s_axi_wstrb
	wire         mm_interconnect_0_axi_adrv9001_s_axi_wready;             // axi_adrv9001:s_axi_wready -> mm_interconnect_0:axi_adrv9001_s_axi_wready
	wire         mm_interconnect_0_axi_adrv9001_s_axi_awready;            // axi_adrv9001:s_axi_awready -> mm_interconnect_0:axi_adrv9001_s_axi_awready
	wire         mm_interconnect_0_axi_adrv9001_s_axi_rready;             // mm_interconnect_0:axi_adrv9001_s_axi_rready -> axi_adrv9001:s_axi_rready
	wire         mm_interconnect_0_axi_adrv9001_s_axi_bready;             // mm_interconnect_0:axi_adrv9001_s_axi_bready -> axi_adrv9001:s_axi_bready
	wire         mm_interconnect_0_axi_adrv9001_s_axi_wvalid;             // mm_interconnect_0:axi_adrv9001_s_axi_wvalid -> axi_adrv9001:s_axi_wvalid
	wire  [15:0] mm_interconnect_0_axi_adrv9001_s_axi_araddr;             // mm_interconnect_0:axi_adrv9001_s_axi_araddr -> axi_adrv9001:s_axi_araddr
	wire   [2:0] mm_interconnect_0_axi_adrv9001_s_axi_arprot;             // mm_interconnect_0:axi_adrv9001_s_axi_arprot -> axi_adrv9001:s_axi_arprot
	wire   [1:0] mm_interconnect_0_axi_adrv9001_s_axi_rresp;              // axi_adrv9001:s_axi_rresp -> mm_interconnect_0:axi_adrv9001_s_axi_rresp
	wire   [2:0] mm_interconnect_0_axi_adrv9001_s_axi_awprot;             // mm_interconnect_0:axi_adrv9001_s_axi_awprot -> axi_adrv9001:s_axi_awprot
	wire  [31:0] mm_interconnect_0_axi_adrv9001_s_axi_wdata;              // mm_interconnect_0:axi_adrv9001_s_axi_wdata -> axi_adrv9001:s_axi_wdata
	wire         mm_interconnect_0_axi_adrv9001_s_axi_arvalid;            // mm_interconnect_0:axi_adrv9001_s_axi_arvalid -> axi_adrv9001:s_axi_arvalid
	wire         mm_interconnect_0_axi_adrv9001_s_axi_bvalid;             // axi_adrv9001:s_axi_bvalid -> mm_interconnect_0:axi_adrv9001_s_axi_bvalid
	wire         mm_interconnect_0_axi_adrv9001_s_axi_awvalid;            // mm_interconnect_0:axi_adrv9001_s_axi_awvalid -> axi_adrv9001:s_axi_awvalid
	wire         mm_interconnect_0_axi_adrv9001_s_axi_rvalid;             // axi_adrv9001:s_axi_rvalid -> mm_interconnect_0:axi_adrv9001_s_axi_rvalid
	wire  [10:0] mm_interconnect_0_axi_adc_dma_s_axi_awaddr;              // mm_interconnect_0:axi_adc_dma_s_axi_awaddr -> axi_adc_dma:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_axi_adc_dma_s_axi_bresp;               // axi_adc_dma:s_axi_bresp -> mm_interconnect_0:axi_adc_dma_s_axi_bresp
	wire         mm_interconnect_0_axi_adc_dma_s_axi_arready;             // axi_adc_dma:s_axi_arready -> mm_interconnect_0:axi_adc_dma_s_axi_arready
	wire  [31:0] mm_interconnect_0_axi_adc_dma_s_axi_rdata;               // axi_adc_dma:s_axi_rdata -> mm_interconnect_0:axi_adc_dma_s_axi_rdata
	wire   [3:0] mm_interconnect_0_axi_adc_dma_s_axi_wstrb;               // mm_interconnect_0:axi_adc_dma_s_axi_wstrb -> axi_adc_dma:s_axi_wstrb
	wire         mm_interconnect_0_axi_adc_dma_s_axi_wready;              // axi_adc_dma:s_axi_wready -> mm_interconnect_0:axi_adc_dma_s_axi_wready
	wire         mm_interconnect_0_axi_adc_dma_s_axi_awready;             // axi_adc_dma:s_axi_awready -> mm_interconnect_0:axi_adc_dma_s_axi_awready
	wire         mm_interconnect_0_axi_adc_dma_s_axi_rready;              // mm_interconnect_0:axi_adc_dma_s_axi_rready -> axi_adc_dma:s_axi_rready
	wire         mm_interconnect_0_axi_adc_dma_s_axi_bready;              // mm_interconnect_0:axi_adc_dma_s_axi_bready -> axi_adc_dma:s_axi_bready
	wire         mm_interconnect_0_axi_adc_dma_s_axi_wvalid;              // mm_interconnect_0:axi_adc_dma_s_axi_wvalid -> axi_adc_dma:s_axi_wvalid
	wire  [10:0] mm_interconnect_0_axi_adc_dma_s_axi_araddr;              // mm_interconnect_0:axi_adc_dma_s_axi_araddr -> axi_adc_dma:s_axi_araddr
	wire   [2:0] mm_interconnect_0_axi_adc_dma_s_axi_arprot;              // mm_interconnect_0:axi_adc_dma_s_axi_arprot -> axi_adc_dma:s_axi_arprot
	wire   [1:0] mm_interconnect_0_axi_adc_dma_s_axi_rresp;               // axi_adc_dma:s_axi_rresp -> mm_interconnect_0:axi_adc_dma_s_axi_rresp
	wire   [2:0] mm_interconnect_0_axi_adc_dma_s_axi_awprot;              // mm_interconnect_0:axi_adc_dma_s_axi_awprot -> axi_adc_dma:s_axi_awprot
	wire  [31:0] mm_interconnect_0_axi_adc_dma_s_axi_wdata;               // mm_interconnect_0:axi_adc_dma_s_axi_wdata -> axi_adc_dma:s_axi_wdata
	wire         mm_interconnect_0_axi_adc_dma_s_axi_arvalid;             // mm_interconnect_0:axi_adc_dma_s_axi_arvalid -> axi_adc_dma:s_axi_arvalid
	wire         mm_interconnect_0_axi_adc_dma_s_axi_bvalid;              // axi_adc_dma:s_axi_bvalid -> mm_interconnect_0:axi_adc_dma_s_axi_bvalid
	wire         mm_interconnect_0_axi_adc_dma_s_axi_awvalid;             // mm_interconnect_0:axi_adc_dma_s_axi_awvalid -> axi_adc_dma:s_axi_awvalid
	wire         mm_interconnect_0_axi_adc_dma_s_axi_rvalid;              // axi_adc_dma:s_axi_rvalid -> mm_interconnect_0:axi_adc_dma_s_axi_rvalid
	wire  [10:0] mm_interconnect_0_axi_dac_dma_s_axi_awaddr;              // mm_interconnect_0:axi_dac_dma_s_axi_awaddr -> axi_dac_dma:s_axi_awaddr
	wire   [1:0] mm_interconnect_0_axi_dac_dma_s_axi_bresp;               // axi_dac_dma:s_axi_bresp -> mm_interconnect_0:axi_dac_dma_s_axi_bresp
	wire         mm_interconnect_0_axi_dac_dma_s_axi_arready;             // axi_dac_dma:s_axi_arready -> mm_interconnect_0:axi_dac_dma_s_axi_arready
	wire  [31:0] mm_interconnect_0_axi_dac_dma_s_axi_rdata;               // axi_dac_dma:s_axi_rdata -> mm_interconnect_0:axi_dac_dma_s_axi_rdata
	wire   [3:0] mm_interconnect_0_axi_dac_dma_s_axi_wstrb;               // mm_interconnect_0:axi_dac_dma_s_axi_wstrb -> axi_dac_dma:s_axi_wstrb
	wire         mm_interconnect_0_axi_dac_dma_s_axi_wready;              // axi_dac_dma:s_axi_wready -> mm_interconnect_0:axi_dac_dma_s_axi_wready
	wire         mm_interconnect_0_axi_dac_dma_s_axi_awready;             // axi_dac_dma:s_axi_awready -> mm_interconnect_0:axi_dac_dma_s_axi_awready
	wire         mm_interconnect_0_axi_dac_dma_s_axi_rready;              // mm_interconnect_0:axi_dac_dma_s_axi_rready -> axi_dac_dma:s_axi_rready
	wire         mm_interconnect_0_axi_dac_dma_s_axi_bready;              // mm_interconnect_0:axi_dac_dma_s_axi_bready -> axi_dac_dma:s_axi_bready
	wire         mm_interconnect_0_axi_dac_dma_s_axi_wvalid;              // mm_interconnect_0:axi_dac_dma_s_axi_wvalid -> axi_dac_dma:s_axi_wvalid
	wire  [10:0] mm_interconnect_0_axi_dac_dma_s_axi_araddr;              // mm_interconnect_0:axi_dac_dma_s_axi_araddr -> axi_dac_dma:s_axi_araddr
	wire   [2:0] mm_interconnect_0_axi_dac_dma_s_axi_arprot;              // mm_interconnect_0:axi_dac_dma_s_axi_arprot -> axi_dac_dma:s_axi_arprot
	wire   [1:0] mm_interconnect_0_axi_dac_dma_s_axi_rresp;               // axi_dac_dma:s_axi_rresp -> mm_interconnect_0:axi_dac_dma_s_axi_rresp
	wire   [2:0] mm_interconnect_0_axi_dac_dma_s_axi_awprot;              // mm_interconnect_0:axi_dac_dma_s_axi_awprot -> axi_dac_dma:s_axi_awprot
	wire  [31:0] mm_interconnect_0_axi_dac_dma_s_axi_wdata;               // mm_interconnect_0:axi_dac_dma_s_axi_wdata -> axi_dac_dma:s_axi_wdata
	wire         mm_interconnect_0_axi_dac_dma_s_axi_arvalid;             // mm_interconnect_0:axi_dac_dma_s_axi_arvalid -> axi_dac_dma:s_axi_arvalid
	wire         mm_interconnect_0_axi_dac_dma_s_axi_bvalid;              // axi_dac_dma:s_axi_bvalid -> mm_interconnect_0:axi_dac_dma_s_axi_bvalid
	wire         mm_interconnect_0_axi_dac_dma_s_axi_awvalid;             // mm_interconnect_0:axi_dac_dma_s_axi_awvalid -> axi_dac_dma:s_axi_awvalid
	wire         mm_interconnect_0_axi_dac_dma_s_axi_rvalid;              // axi_dac_dma:s_axi_rvalid -> mm_interconnect_0:axi_dac_dma_s_axi_rvalid
	wire         mm_interconnect_0_spi_0_spi_control_port_chipselect;     // mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_readdata;       // spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_spi_0_spi_control_port_address;        // mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	wire         mm_interconnect_0_spi_0_spi_control_port_read;           // mm_interconnect_0:spi_0_spi_control_port_read -> spi_0:read_n
	wire         mm_interconnect_0_spi_0_spi_control_port_write;          // mm_interconnect_0:spi_0_spi_control_port_write -> spi_0:write_n
	wire  [15:0] mm_interconnect_0_spi_0_spi_control_port_writedata;      // mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	wire   [1:0] axi_adc_dma_m_dest_axi_awburst;                          // axi_adc_dma:m_dest_axi_awburst -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awburst
	wire   [3:0] axi_adc_dma_m_dest_axi_arlen;                            // axi_adc_dma:m_dest_axi_arlen -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arlen
	wire   [7:0] axi_adc_dma_m_dest_axi_wstrb;                            // axi_adc_dma:m_dest_axi_wstrb -> mm_interconnect_1:axi_adc_dma_m_dest_axi_wstrb
	wire         axi_adc_dma_m_dest_axi_wready;                           // mm_interconnect_1:axi_adc_dma_m_dest_axi_wready -> axi_adc_dma:m_dest_axi_wready
	wire         axi_adc_dma_m_dest_axi_rid;                              // mm_interconnect_1:axi_adc_dma_m_dest_axi_rid -> axi_adc_dma:m_dest_axi_rid
	wire         axi_adc_dma_m_dest_axi_rready;                           // axi_adc_dma:m_dest_axi_rready -> mm_interconnect_1:axi_adc_dma_m_dest_axi_rready
	wire   [3:0] axi_adc_dma_m_dest_axi_awlen;                            // axi_adc_dma:m_dest_axi_awlen -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awlen
	wire         axi_adc_dma_m_dest_axi_wid;                              // axi_adc_dma:m_dest_axi_wid -> mm_interconnect_1:axi_adc_dma_m_dest_axi_wid
	wire   [3:0] axi_adc_dma_m_dest_axi_arcache;                          // axi_adc_dma:m_dest_axi_arcache -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arcache
	wire         axi_adc_dma_m_dest_axi_wvalid;                           // axi_adc_dma:m_dest_axi_wvalid -> mm_interconnect_1:axi_adc_dma_m_dest_axi_wvalid
	wire  [31:0] axi_adc_dma_m_dest_axi_araddr;                           // axi_adc_dma:m_dest_axi_araddr -> mm_interconnect_1:axi_adc_dma_m_dest_axi_araddr
	wire   [2:0] axi_adc_dma_m_dest_axi_arprot;                           // axi_adc_dma:m_dest_axi_arprot -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arprot
	wire  [63:0] axi_adc_dma_m_dest_axi_wdata;                            // axi_adc_dma:m_dest_axi_wdata -> mm_interconnect_1:axi_adc_dma_m_dest_axi_wdata
	wire         axi_adc_dma_m_dest_axi_arvalid;                          // axi_adc_dma:m_dest_axi_arvalid -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arvalid
	wire   [2:0] axi_adc_dma_m_dest_axi_awprot;                           // axi_adc_dma:m_dest_axi_awprot -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awprot
	wire   [3:0] axi_adc_dma_m_dest_axi_awcache;                          // axi_adc_dma:m_dest_axi_awcache -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awcache
	wire         axi_adc_dma_m_dest_axi_arid;                             // axi_adc_dma:m_dest_axi_arid -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arid
	wire   [1:0] axi_adc_dma_m_dest_axi_arlock;                           // axi_adc_dma:m_dest_axi_arlock -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arlock
	wire   [1:0] axi_adc_dma_m_dest_axi_awlock;                           // axi_adc_dma:m_dest_axi_awlock -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awlock
	wire  [31:0] axi_adc_dma_m_dest_axi_awaddr;                           // axi_adc_dma:m_dest_axi_awaddr -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awaddr
	wire   [1:0] axi_adc_dma_m_dest_axi_bresp;                            // mm_interconnect_1:axi_adc_dma_m_dest_axi_bresp -> axi_adc_dma:m_dest_axi_bresp
	wire         axi_adc_dma_m_dest_axi_arready;                          // mm_interconnect_1:axi_adc_dma_m_dest_axi_arready -> axi_adc_dma:m_dest_axi_arready
	wire  [63:0] axi_adc_dma_m_dest_axi_rdata;                            // mm_interconnect_1:axi_adc_dma_m_dest_axi_rdata -> axi_adc_dma:m_dest_axi_rdata
	wire         axi_adc_dma_m_dest_axi_awready;                          // mm_interconnect_1:axi_adc_dma_m_dest_axi_awready -> axi_adc_dma:m_dest_axi_awready
	wire   [1:0] axi_adc_dma_m_dest_axi_arburst;                          // axi_adc_dma:m_dest_axi_arburst -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arburst
	wire   [2:0] axi_adc_dma_m_dest_axi_arsize;                           // axi_adc_dma:m_dest_axi_arsize -> mm_interconnect_1:axi_adc_dma_m_dest_axi_arsize
	wire         axi_adc_dma_m_dest_axi_bready;                           // axi_adc_dma:m_dest_axi_bready -> mm_interconnect_1:axi_adc_dma_m_dest_axi_bready
	wire         axi_adc_dma_m_dest_axi_rlast;                            // mm_interconnect_1:axi_adc_dma_m_dest_axi_rlast -> axi_adc_dma:m_dest_axi_rlast
	wire         axi_adc_dma_m_dest_axi_wlast;                            // axi_adc_dma:m_dest_axi_wlast -> mm_interconnect_1:axi_adc_dma_m_dest_axi_wlast
	wire   [1:0] axi_adc_dma_m_dest_axi_rresp;                            // mm_interconnect_1:axi_adc_dma_m_dest_axi_rresp -> axi_adc_dma:m_dest_axi_rresp
	wire         axi_adc_dma_m_dest_axi_awid;                             // axi_adc_dma:m_dest_axi_awid -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awid
	wire         axi_adc_dma_m_dest_axi_bid;                              // mm_interconnect_1:axi_adc_dma_m_dest_axi_bid -> axi_adc_dma:m_dest_axi_bid
	wire         axi_adc_dma_m_dest_axi_bvalid;                           // mm_interconnect_1:axi_adc_dma_m_dest_axi_bvalid -> axi_adc_dma:m_dest_axi_bvalid
	wire         axi_adc_dma_m_dest_axi_awvalid;                          // axi_adc_dma:m_dest_axi_awvalid -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awvalid
	wire         axi_adc_dma_m_dest_axi_rvalid;                           // mm_interconnect_1:axi_adc_dma_m_dest_axi_rvalid -> axi_adc_dma:m_dest_axi_rvalid
	wire   [2:0] axi_adc_dma_m_dest_axi_awsize;                           // axi_adc_dma:m_dest_axi_awsize -> mm_interconnect_1:axi_adc_dma_m_dest_axi_awsize
	wire   [1:0] hdmi_dmac_0_m_src_axi_awburst;                           // hdmi_dmac_0:m_src_axi_awburst -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awburst
	wire   [3:0] hdmi_dmac_0_m_src_axi_arlen;                             // hdmi_dmac_0:m_src_axi_arlen -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arlen
	wire   [7:0] hdmi_dmac_0_m_src_axi_wstrb;                             // hdmi_dmac_0:m_src_axi_wstrb -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_wstrb
	wire         hdmi_dmac_0_m_src_axi_wready;                            // mm_interconnect_1:hdmi_dmac_0_m_src_axi_wready -> hdmi_dmac_0:m_src_axi_wready
	wire         hdmi_dmac_0_m_src_axi_rid;                               // mm_interconnect_1:hdmi_dmac_0_m_src_axi_rid -> hdmi_dmac_0:m_src_axi_rid
	wire         hdmi_dmac_0_m_src_axi_rready;                            // hdmi_dmac_0:m_src_axi_rready -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_rready
	wire   [3:0] hdmi_dmac_0_m_src_axi_awlen;                             // hdmi_dmac_0:m_src_axi_awlen -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awlen
	wire         hdmi_dmac_0_m_src_axi_wid;                               // hdmi_dmac_0:m_src_axi_wid -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_wid
	wire   [3:0] hdmi_dmac_0_m_src_axi_arcache;                           // hdmi_dmac_0:m_src_axi_arcache -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arcache
	wire         hdmi_dmac_0_m_src_axi_wvalid;                            // hdmi_dmac_0:m_src_axi_wvalid -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_wvalid
	wire  [31:0] hdmi_dmac_0_m_src_axi_araddr;                            // hdmi_dmac_0:m_src_axi_araddr -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_araddr
	wire   [2:0] hdmi_dmac_0_m_src_axi_arprot;                            // hdmi_dmac_0:m_src_axi_arprot -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arprot
	wire  [63:0] hdmi_dmac_0_m_src_axi_wdata;                             // hdmi_dmac_0:m_src_axi_wdata -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_wdata
	wire         hdmi_dmac_0_m_src_axi_arvalid;                           // hdmi_dmac_0:m_src_axi_arvalid -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arvalid
	wire   [2:0] hdmi_dmac_0_m_src_axi_awprot;                            // hdmi_dmac_0:m_src_axi_awprot -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awprot
	wire   [3:0] hdmi_dmac_0_m_src_axi_awcache;                           // hdmi_dmac_0:m_src_axi_awcache -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awcache
	wire         hdmi_dmac_0_m_src_axi_arid;                              // hdmi_dmac_0:m_src_axi_arid -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arid
	wire   [1:0] hdmi_dmac_0_m_src_axi_arlock;                            // hdmi_dmac_0:m_src_axi_arlock -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arlock
	wire   [1:0] hdmi_dmac_0_m_src_axi_awlock;                            // hdmi_dmac_0:m_src_axi_awlock -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awlock
	wire  [31:0] hdmi_dmac_0_m_src_axi_awaddr;                            // hdmi_dmac_0:m_src_axi_awaddr -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awaddr
	wire   [1:0] hdmi_dmac_0_m_src_axi_bresp;                             // mm_interconnect_1:hdmi_dmac_0_m_src_axi_bresp -> hdmi_dmac_0:m_src_axi_bresp
	wire         hdmi_dmac_0_m_src_axi_arready;                           // mm_interconnect_1:hdmi_dmac_0_m_src_axi_arready -> hdmi_dmac_0:m_src_axi_arready
	wire  [63:0] hdmi_dmac_0_m_src_axi_rdata;                             // mm_interconnect_1:hdmi_dmac_0_m_src_axi_rdata -> hdmi_dmac_0:m_src_axi_rdata
	wire         hdmi_dmac_0_m_src_axi_awready;                           // mm_interconnect_1:hdmi_dmac_0_m_src_axi_awready -> hdmi_dmac_0:m_src_axi_awready
	wire   [1:0] hdmi_dmac_0_m_src_axi_arburst;                           // hdmi_dmac_0:m_src_axi_arburst -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arburst
	wire   [2:0] hdmi_dmac_0_m_src_axi_arsize;                            // hdmi_dmac_0:m_src_axi_arsize -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_arsize
	wire         hdmi_dmac_0_m_src_axi_bready;                            // hdmi_dmac_0:m_src_axi_bready -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_bready
	wire         hdmi_dmac_0_m_src_axi_rlast;                             // mm_interconnect_1:hdmi_dmac_0_m_src_axi_rlast -> hdmi_dmac_0:m_src_axi_rlast
	wire         hdmi_dmac_0_m_src_axi_wlast;                             // hdmi_dmac_0:m_src_axi_wlast -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_wlast
	wire   [1:0] hdmi_dmac_0_m_src_axi_rresp;                             // mm_interconnect_1:hdmi_dmac_0_m_src_axi_rresp -> hdmi_dmac_0:m_src_axi_rresp
	wire         hdmi_dmac_0_m_src_axi_awid;                              // hdmi_dmac_0:m_src_axi_awid -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awid
	wire         hdmi_dmac_0_m_src_axi_bid;                               // mm_interconnect_1:hdmi_dmac_0_m_src_axi_bid -> hdmi_dmac_0:m_src_axi_bid
	wire         hdmi_dmac_0_m_src_axi_bvalid;                            // mm_interconnect_1:hdmi_dmac_0_m_src_axi_bvalid -> hdmi_dmac_0:m_src_axi_bvalid
	wire         hdmi_dmac_0_m_src_axi_awvalid;                           // hdmi_dmac_0:m_src_axi_awvalid -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awvalid
	wire         hdmi_dmac_0_m_src_axi_rvalid;                            // mm_interconnect_1:hdmi_dmac_0_m_src_axi_rvalid -> hdmi_dmac_0:m_src_axi_rvalid
	wire   [2:0] hdmi_dmac_0_m_src_axi_awsize;                            // hdmi_dmac_0:m_src_axi_awsize -> mm_interconnect_1:hdmi_dmac_0_m_src_axi_awsize
	wire   [1:0] axi_dac_dma_m_src_axi_awburst;                           // axi_dac_dma:m_src_axi_awburst -> mm_interconnect_1:axi_dac_dma_m_src_axi_awburst
	wire   [3:0] axi_dac_dma_m_src_axi_arlen;                             // axi_dac_dma:m_src_axi_arlen -> mm_interconnect_1:axi_dac_dma_m_src_axi_arlen
	wire   [7:0] axi_dac_dma_m_src_axi_wstrb;                             // axi_dac_dma:m_src_axi_wstrb -> mm_interconnect_1:axi_dac_dma_m_src_axi_wstrb
	wire         axi_dac_dma_m_src_axi_wready;                            // mm_interconnect_1:axi_dac_dma_m_src_axi_wready -> axi_dac_dma:m_src_axi_wready
	wire         axi_dac_dma_m_src_axi_rid;                               // mm_interconnect_1:axi_dac_dma_m_src_axi_rid -> axi_dac_dma:m_src_axi_rid
	wire         axi_dac_dma_m_src_axi_rready;                            // axi_dac_dma:m_src_axi_rready -> mm_interconnect_1:axi_dac_dma_m_src_axi_rready
	wire   [3:0] axi_dac_dma_m_src_axi_awlen;                             // axi_dac_dma:m_src_axi_awlen -> mm_interconnect_1:axi_dac_dma_m_src_axi_awlen
	wire         axi_dac_dma_m_src_axi_wid;                               // axi_dac_dma:m_src_axi_wid -> mm_interconnect_1:axi_dac_dma_m_src_axi_wid
	wire   [3:0] axi_dac_dma_m_src_axi_arcache;                           // axi_dac_dma:m_src_axi_arcache -> mm_interconnect_1:axi_dac_dma_m_src_axi_arcache
	wire         axi_dac_dma_m_src_axi_wvalid;                            // axi_dac_dma:m_src_axi_wvalid -> mm_interconnect_1:axi_dac_dma_m_src_axi_wvalid
	wire  [31:0] axi_dac_dma_m_src_axi_araddr;                            // axi_dac_dma:m_src_axi_araddr -> mm_interconnect_1:axi_dac_dma_m_src_axi_araddr
	wire   [2:0] axi_dac_dma_m_src_axi_arprot;                            // axi_dac_dma:m_src_axi_arprot -> mm_interconnect_1:axi_dac_dma_m_src_axi_arprot
	wire  [63:0] axi_dac_dma_m_src_axi_wdata;                             // axi_dac_dma:m_src_axi_wdata -> mm_interconnect_1:axi_dac_dma_m_src_axi_wdata
	wire         axi_dac_dma_m_src_axi_arvalid;                           // axi_dac_dma:m_src_axi_arvalid -> mm_interconnect_1:axi_dac_dma_m_src_axi_arvalid
	wire   [2:0] axi_dac_dma_m_src_axi_awprot;                            // axi_dac_dma:m_src_axi_awprot -> mm_interconnect_1:axi_dac_dma_m_src_axi_awprot
	wire   [3:0] axi_dac_dma_m_src_axi_awcache;                           // axi_dac_dma:m_src_axi_awcache -> mm_interconnect_1:axi_dac_dma_m_src_axi_awcache
	wire         axi_dac_dma_m_src_axi_arid;                              // axi_dac_dma:m_src_axi_arid -> mm_interconnect_1:axi_dac_dma_m_src_axi_arid
	wire   [1:0] axi_dac_dma_m_src_axi_arlock;                            // axi_dac_dma:m_src_axi_arlock -> mm_interconnect_1:axi_dac_dma_m_src_axi_arlock
	wire   [1:0] axi_dac_dma_m_src_axi_awlock;                            // axi_dac_dma:m_src_axi_awlock -> mm_interconnect_1:axi_dac_dma_m_src_axi_awlock
	wire  [31:0] axi_dac_dma_m_src_axi_awaddr;                            // axi_dac_dma:m_src_axi_awaddr -> mm_interconnect_1:axi_dac_dma_m_src_axi_awaddr
	wire   [1:0] axi_dac_dma_m_src_axi_bresp;                             // mm_interconnect_1:axi_dac_dma_m_src_axi_bresp -> axi_dac_dma:m_src_axi_bresp
	wire         axi_dac_dma_m_src_axi_arready;                           // mm_interconnect_1:axi_dac_dma_m_src_axi_arready -> axi_dac_dma:m_src_axi_arready
	wire  [63:0] axi_dac_dma_m_src_axi_rdata;                             // mm_interconnect_1:axi_dac_dma_m_src_axi_rdata -> axi_dac_dma:m_src_axi_rdata
	wire         axi_dac_dma_m_src_axi_awready;                           // mm_interconnect_1:axi_dac_dma_m_src_axi_awready -> axi_dac_dma:m_src_axi_awready
	wire   [1:0] axi_dac_dma_m_src_axi_arburst;                           // axi_dac_dma:m_src_axi_arburst -> mm_interconnect_1:axi_dac_dma_m_src_axi_arburst
	wire   [2:0] axi_dac_dma_m_src_axi_arsize;                            // axi_dac_dma:m_src_axi_arsize -> mm_interconnect_1:axi_dac_dma_m_src_axi_arsize
	wire         axi_dac_dma_m_src_axi_bready;                            // axi_dac_dma:m_src_axi_bready -> mm_interconnect_1:axi_dac_dma_m_src_axi_bready
	wire         axi_dac_dma_m_src_axi_rlast;                             // mm_interconnect_1:axi_dac_dma_m_src_axi_rlast -> axi_dac_dma:m_src_axi_rlast
	wire         axi_dac_dma_m_src_axi_wlast;                             // axi_dac_dma:m_src_axi_wlast -> mm_interconnect_1:axi_dac_dma_m_src_axi_wlast
	wire   [1:0] axi_dac_dma_m_src_axi_rresp;                             // mm_interconnect_1:axi_dac_dma_m_src_axi_rresp -> axi_dac_dma:m_src_axi_rresp
	wire         axi_dac_dma_m_src_axi_awid;                              // axi_dac_dma:m_src_axi_awid -> mm_interconnect_1:axi_dac_dma_m_src_axi_awid
	wire         axi_dac_dma_m_src_axi_bid;                               // mm_interconnect_1:axi_dac_dma_m_src_axi_bid -> axi_dac_dma:m_src_axi_bid
	wire         axi_dac_dma_m_src_axi_bvalid;                            // mm_interconnect_1:axi_dac_dma_m_src_axi_bvalid -> axi_dac_dma:m_src_axi_bvalid
	wire         axi_dac_dma_m_src_axi_awvalid;                           // axi_dac_dma:m_src_axi_awvalid -> mm_interconnect_1:axi_dac_dma_m_src_axi_awvalid
	wire         axi_dac_dma_m_src_axi_rvalid;                            // mm_interconnect_1:axi_dac_dma_m_src_axi_rvalid -> axi_dac_dma:m_src_axi_rvalid
	wire   [2:0] axi_dac_dma_m_src_axi_awsize;                            // axi_dac_dma:m_src_axi_awsize -> mm_interconnect_1:axi_dac_dma_m_src_axi_awsize
	wire  [63:0] mm_interconnect_1_sys_hps_f2h_sdram0_data_readdata;      // sys_hps:f2h_sdram0_READDATA -> mm_interconnect_1:sys_hps_f2h_sdram0_data_readdata
	wire         mm_interconnect_1_sys_hps_f2h_sdram0_data_waitrequest;   // sys_hps:f2h_sdram0_WAITREQUEST -> mm_interconnect_1:sys_hps_f2h_sdram0_data_waitrequest
	wire  [28:0] mm_interconnect_1_sys_hps_f2h_sdram0_data_address;       // mm_interconnect_1:sys_hps_f2h_sdram0_data_address -> sys_hps:f2h_sdram0_ADDRESS
	wire         mm_interconnect_1_sys_hps_f2h_sdram0_data_read;          // mm_interconnect_1:sys_hps_f2h_sdram0_data_read -> sys_hps:f2h_sdram0_READ
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram0_data_byteenable;    // mm_interconnect_1:sys_hps_f2h_sdram0_data_byteenable -> sys_hps:f2h_sdram0_BYTEENABLE
	wire         mm_interconnect_1_sys_hps_f2h_sdram0_data_readdatavalid; // sys_hps:f2h_sdram0_READDATAVALID -> mm_interconnect_1:sys_hps_f2h_sdram0_data_readdatavalid
	wire         mm_interconnect_1_sys_hps_f2h_sdram0_data_write;         // mm_interconnect_1:sys_hps_f2h_sdram0_data_write -> sys_hps:f2h_sdram0_WRITE
	wire  [63:0] mm_interconnect_1_sys_hps_f2h_sdram0_data_writedata;     // mm_interconnect_1:sys_hps_f2h_sdram0_data_writedata -> sys_hps:f2h_sdram0_WRITEDATA
	wire   [7:0] mm_interconnect_1_sys_hps_f2h_sdram0_data_burstcount;    // mm_interconnect_1:sys_hps_f2h_sdram0_data_burstcount -> sys_hps:f2h_sdram0_BURSTCOUNT
	wire         irq_mapper_receiver0_irq;                                // hdmi_dmac_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                // axi_adc_dma:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                // axi_dac_dma:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                // sys_gpio_bd:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                // sys_gpio_in:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                // spi_0:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                // avl_adrv9001_gpio:irq -> irq_mapper:receiver6_irq
	wire  [31:0] sys_hps_f2h_irq0_irq;                                    // irq_mapper:sender_irq -> sys_hps:f2h_irq_p0
	wire  [31:0] sys_hps_f2h_irq1_irq;                                    // irq_mapper_001:sender_irq -> sys_hps:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [avl_adrv9001_gpio:reset_n, axi_adc_dma:m_dest_axi_aresetn, axi_adc_dma:s_axi_aresetn, axi_adrv9001:s_axi_aresetn, axi_dac_dma:m_src_axi_aresetn, axi_dac_dma:s_axi_aresetn, axi_hdmi_tx_0:s_axi_aresetn, hdmi_dmac_0:m_src_axi_aresetn, hdmi_dmac_0:s_axi_aresetn, mm_interconnect_0:sys_id_reset_reset_bridge_in_reset_reset, mm_interconnect_1:axi_adc_dma_m_dest_axi_reset_reset_bridge_in_reset_reset, spi_0:reset_n, sys_gpio_bd:reset_n, sys_gpio_in:reset_n, sys_gpio_out:reset_n, sys_id:reset_n, util_adc_pack:reset, util_adc_wfifo:dout_rstn, util_dac_rfifo:din_rstn, util_dac_upack:reset]
	wire         rst_controller_001_reset_out_reset;                      // rst_controller_001:reset_out -> [mm_interconnect_0:sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sys_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset]
	wire   [0:0] util_dac_upack_fifo_rd_valid;                            // port fragment
	wire  [63:0] util_dac_upack_fifo_rd_data;                             // port fragment

	system_bd_avl_adrv9001_gpio avl_adrv9001_gpio (
		.clk        (sys_hps_h2f_user1_clock_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address    (mm_interconnect_0_avl_adrv9001_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_avl_adrv9001_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_avl_adrv9001_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_avl_adrv9001_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_avl_adrv9001_gpio_s1_readdata),   //                    .readdata
		.bidir_port (adrv9001_gpio_export),                              // external_connection.export
		.irq        (irq_mapper_receiver6_irq)                           //                 irq.irq
	);

	axi_dmac #(
		.ID                    (0),
		.DMA_LENGTH_WIDTH      (24),
		.FIFO_SIZE             (4),
		.MAX_BYTES_PER_BURST   (128),
		.DMA_TYPE_SRC          (2),
		.DMA_AXI_PROTOCOL_SRC  (1),
		.DMA_DATA_WIDTH_SRC    (64),
		.AXI_SLICE_SRC         (0),
		.DMA_TYPE_DEST         (0),
		.DMA_AXI_PROTOCOL_DEST (1),
		.DMA_DATA_WIDTH_DEST   (64),
		.AXI_SLICE_DEST        (0),
		.CYCLIC                (0),
		.DMA_2D_TRANSFER       (0),
		.SYNC_TRANSFER_START   (1),
		.ASYNC_CLK_REQ_SRC     (0),
		.ASYNC_CLK_SRC_DEST    (0),
		.ASYNC_CLK_DEST_REQ    (0),
		.ENABLE_DIAGNOSTICS_IF (0),
		.DMA_AXIS_ID_W         (8),
		.DMA_AXIS_DEST_W       (4)
	) axi_adc_dma (
		.s_axi_aclk             (sys_hps_h2f_user1_clock_clk),                                          //         s_axi_clock.clk
		.s_axi_aresetn          (~rst_controller_reset_out_reset),                                      //         s_axi_reset.reset_n
		.s_axi_awvalid          (mm_interconnect_0_axi_adc_dma_s_axi_awvalid),                          //               s_axi.awvalid
		.s_axi_awaddr           (mm_interconnect_0_axi_adc_dma_s_axi_awaddr),                           //                    .awaddr
		.s_axi_awprot           (mm_interconnect_0_axi_adc_dma_s_axi_awprot),                           //                    .awprot
		.s_axi_awready          (mm_interconnect_0_axi_adc_dma_s_axi_awready),                          //                    .awready
		.s_axi_wvalid           (mm_interconnect_0_axi_adc_dma_s_axi_wvalid),                           //                    .wvalid
		.s_axi_wdata            (mm_interconnect_0_axi_adc_dma_s_axi_wdata),                            //                    .wdata
		.s_axi_wstrb            (mm_interconnect_0_axi_adc_dma_s_axi_wstrb),                            //                    .wstrb
		.s_axi_wready           (mm_interconnect_0_axi_adc_dma_s_axi_wready),                           //                    .wready
		.s_axi_bvalid           (mm_interconnect_0_axi_adc_dma_s_axi_bvalid),                           //                    .bvalid
		.s_axi_bresp            (mm_interconnect_0_axi_adc_dma_s_axi_bresp),                            //                    .bresp
		.s_axi_bready           (mm_interconnect_0_axi_adc_dma_s_axi_bready),                           //                    .bready
		.s_axi_arvalid          (mm_interconnect_0_axi_adc_dma_s_axi_arvalid),                          //                    .arvalid
		.s_axi_araddr           (mm_interconnect_0_axi_adc_dma_s_axi_araddr),                           //                    .araddr
		.s_axi_arprot           (mm_interconnect_0_axi_adc_dma_s_axi_arprot),                           //                    .arprot
		.s_axi_arready          (mm_interconnect_0_axi_adc_dma_s_axi_arready),                          //                    .arready
		.s_axi_rvalid           (mm_interconnect_0_axi_adc_dma_s_axi_rvalid),                           //                    .rvalid
		.s_axi_rresp            (mm_interconnect_0_axi_adc_dma_s_axi_rresp),                            //                    .rresp
		.s_axi_rdata            (mm_interconnect_0_axi_adc_dma_s_axi_rdata),                            //                    .rdata
		.s_axi_rready           (mm_interconnect_0_axi_adc_dma_s_axi_rready),                           //                    .rready
		.irq                    (irq_mapper_receiver1_irq),                                             //    interrupt_sender.irq
		.m_dest_axi_aclk        (sys_hps_h2f_user1_clock_clk),                                          //    m_dest_axi_clock.clk
		.m_dest_axi_aresetn     (~rst_controller_reset_out_reset),                                      //    m_dest_axi_reset.reset_n
		.fifo_wr_clk            (sys_hps_h2f_user1_clock_clk),                                          //      if_fifo_wr_clk.clk
		.fifo_wr_en             (util_adc_pack_if_packed_fifo_wr_en_valid),                             //       if_fifo_wr_en.valid
		.fifo_wr_din            (util_adc_pack_if_packed_fifo_wr_data_data),                            //      if_fifo_wr_din.data
		.fifo_wr_overflow       (axi_adc_dma_if_fifo_wr_overflow_ovf),                                  // if_fifo_wr_overflow.ovf
		.fifo_wr_sync           (util_adc_pack_if_packed_fifo_wr_sync_sync),                            //     if_fifo_wr_sync.sync
		.fifo_wr_xfer_req       (),                                                                     // if_fifo_wr_xfer_req.xfer_req
		.m_dest_axi_awvalid     (axi_adc_dma_m_dest_axi_awvalid),                                       //          m_dest_axi.awvalid
		.m_dest_axi_awaddr      (axi_adc_dma_m_dest_axi_awaddr),                                        //                    .awaddr
		.m_dest_axi_awready     (axi_adc_dma_m_dest_axi_awready),                                       //                    .awready
		.m_dest_axi_wvalid      (axi_adc_dma_m_dest_axi_wvalid),                                        //                    .wvalid
		.m_dest_axi_wdata       (axi_adc_dma_m_dest_axi_wdata),                                         //                    .wdata
		.m_dest_axi_wstrb       (axi_adc_dma_m_dest_axi_wstrb),                                         //                    .wstrb
		.m_dest_axi_wready      (axi_adc_dma_m_dest_axi_wready),                                        //                    .wready
		.m_dest_axi_bvalid      (axi_adc_dma_m_dest_axi_bvalid),                                        //                    .bvalid
		.m_dest_axi_bresp       (axi_adc_dma_m_dest_axi_bresp),                                         //                    .bresp
		.m_dest_axi_bready      (axi_adc_dma_m_dest_axi_bready),                                        //                    .bready
		.m_dest_axi_arvalid     (axi_adc_dma_m_dest_axi_arvalid),                                       //                    .arvalid
		.m_dest_axi_araddr      (axi_adc_dma_m_dest_axi_araddr),                                        //                    .araddr
		.m_dest_axi_arready     (axi_adc_dma_m_dest_axi_arready),                                       //                    .arready
		.m_dest_axi_rvalid      (axi_adc_dma_m_dest_axi_rvalid),                                        //                    .rvalid
		.m_dest_axi_rresp       (axi_adc_dma_m_dest_axi_rresp),                                         //                    .rresp
		.m_dest_axi_rdata       (axi_adc_dma_m_dest_axi_rdata),                                         //                    .rdata
		.m_dest_axi_rready      (axi_adc_dma_m_dest_axi_rready),                                        //                    .rready
		.m_dest_axi_awlen       (axi_adc_dma_m_dest_axi_awlen),                                         //                    .awlen
		.m_dest_axi_awsize      (axi_adc_dma_m_dest_axi_awsize),                                        //                    .awsize
		.m_dest_axi_awburst     (axi_adc_dma_m_dest_axi_awburst),                                       //                    .awburst
		.m_dest_axi_awcache     (axi_adc_dma_m_dest_axi_awcache),                                       //                    .awcache
		.m_dest_axi_awprot      (axi_adc_dma_m_dest_axi_awprot),                                        //                    .awprot
		.m_dest_axi_wlast       (axi_adc_dma_m_dest_axi_wlast),                                         //                    .wlast
		.m_dest_axi_arlen       (axi_adc_dma_m_dest_axi_arlen),                                         //                    .arlen
		.m_dest_axi_arsize      (axi_adc_dma_m_dest_axi_arsize),                                        //                    .arsize
		.m_dest_axi_arburst     (axi_adc_dma_m_dest_axi_arburst),                                       //                    .arburst
		.m_dest_axi_arcache     (axi_adc_dma_m_dest_axi_arcache),                                       //                    .arcache
		.m_dest_axi_arprot      (axi_adc_dma_m_dest_axi_arprot),                                        //                    .arprot
		.m_dest_axi_awid        (axi_adc_dma_m_dest_axi_awid),                                          //                    .awid
		.m_dest_axi_awlock      (axi_adc_dma_m_dest_axi_awlock),                                        //                    .awlock
		.m_dest_axi_wid         (axi_adc_dma_m_dest_axi_wid),                                           //                    .wid
		.m_dest_axi_arid        (axi_adc_dma_m_dest_axi_arid),                                          //                    .arid
		.m_dest_axi_arlock      (axi_adc_dma_m_dest_axi_arlock),                                        //                    .arlock
		.m_dest_axi_rid         (axi_adc_dma_m_dest_axi_rid),                                           //                    .rid
		.m_dest_axi_bid         (axi_adc_dma_m_dest_axi_bid),                                           //                    .bid
		.m_dest_axi_rlast       (axi_adc_dma_m_dest_axi_rlast),                                         //                    .rlast
		.m_src_axi_aclk         (1'b0),                                                                 //         (terminated)
		.m_src_axi_aresetn      (1'b1),                                                                 //         (terminated)
		.m_axis_aclk            (1'b0),                                                                 //         (terminated)
		.m_axis_xfer_req        (),                                                                     //         (terminated)
		.m_axis_valid           (),                                                                     //         (terminated)
		.m_axis_last            (),                                                                     //         (terminated)
		.m_axis_ready           (1'b0),                                                                 //         (terminated)
		.m_axis_data            (),                                                                     //         (terminated)
		.m_axis_user            (),                                                                     //         (terminated)
		.m_axis_id              (),                                                                     //         (terminated)
		.m_axis_dest            (),                                                                     //         (terminated)
		.m_axis_strb            (),                                                                     //         (terminated)
		.m_axis_keep            (),                                                                     //         (terminated)
		.s_axis_aclk            (1'b0),                                                                 //         (terminated)
		.s_axis_xfer_req        (),                                                                     //         (terminated)
		.s_axis_valid           (1'b0),                                                                 //         (terminated)
		.s_axis_last            (1'b0),                                                                 //         (terminated)
		.s_axis_ready           (),                                                                     //         (terminated)
		.s_axis_data            (64'b0000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.s_axis_user            (1'b0),                                                                 //         (terminated)
		.s_axis_id              (8'b00000000),                                                          //         (terminated)
		.s_axis_dest            (4'b0000),                                                              //         (terminated)
		.s_axis_strb            (8'b00000000),                                                          //         (terminated)
		.s_axis_keep            (8'b00000000),                                                          //         (terminated)
		.fifo_rd_clk            (1'b0),                                                                 //         (terminated)
		.fifo_rd_en             (1'b0),                                                                 //         (terminated)
		.fifo_rd_valid          (),                                                                     //         (terminated)
		.fifo_rd_dout           (),                                                                     //         (terminated)
		.fifo_rd_underflow      (),                                                                     //         (terminated)
		.fifo_rd_xfer_req       (),                                                                     //         (terminated)
		.dest_diag_level_bursts (),                                                                     //         (terminated)
		.m_src_axi_awvalid      (),                                                                     //         (terminated)
		.m_src_axi_awaddr       (),                                                                     //         (terminated)
		.m_src_axi_awready      (1'b0),                                                                 //         (terminated)
		.m_src_axi_wvalid       (),                                                                     //         (terminated)
		.m_src_axi_wdata        (),                                                                     //         (terminated)
		.m_src_axi_wstrb        (),                                                                     //         (terminated)
		.m_src_axi_wready       (1'b0),                                                                 //         (terminated)
		.m_src_axi_bvalid       (1'b0),                                                                 //         (terminated)
		.m_src_axi_bresp        (2'b00),                                                                //         (terminated)
		.m_src_axi_bready       (),                                                                     //         (terminated)
		.m_src_axi_arvalid      (),                                                                     //         (terminated)
		.m_src_axi_araddr       (),                                                                     //         (terminated)
		.m_src_axi_arready      (1'b0),                                                                 //         (terminated)
		.m_src_axi_rvalid       (1'b0),                                                                 //         (terminated)
		.m_src_axi_rresp        (2'b00),                                                                //         (terminated)
		.m_src_axi_rdata        (64'b0000000000000000000000000000000000000000000000000000000000000000), //         (terminated)
		.m_src_axi_rready       (),                                                                     //         (terminated)
		.m_src_axi_awlen        (),                                                                     //         (terminated)
		.m_src_axi_awsize       (),                                                                     //         (terminated)
		.m_src_axi_awburst      (),                                                                     //         (terminated)
		.m_src_axi_awcache      (),                                                                     //         (terminated)
		.m_src_axi_awprot       (),                                                                     //         (terminated)
		.m_src_axi_wlast        (),                                                                     //         (terminated)
		.m_src_axi_arlen        (),                                                                     //         (terminated)
		.m_src_axi_arsize       (),                                                                     //         (terminated)
		.m_src_axi_arburst      (),                                                                     //         (terminated)
		.m_src_axi_arcache      (),                                                                     //         (terminated)
		.m_src_axi_arprot       (),                                                                     //         (terminated)
		.m_src_axi_awid         (),                                                                     //         (terminated)
		.m_src_axi_awlock       (),                                                                     //         (terminated)
		.m_src_axi_wid          (),                                                                     //         (terminated)
		.m_src_axi_arid         (),                                                                     //         (terminated)
		.m_src_axi_arlock       (),                                                                     //         (terminated)
		.m_src_axi_rid          (1'b0),                                                                 //         (terminated)
		.m_src_axi_bid          (1'b0),                                                                 //         (terminated)
		.m_src_axi_rlast        (1'b0)                                                                  //         (terminated)
	);

	axi_adrv9001 #(
		.ID              (0),
		.CMOS_LVDS_N     (1),
		.IO_DELAY_GROUP  ("dev_if_delay_group"),
		.FPGA_TECHNOLOGY (101),
		.FPGA_FAMILY     (5),
		.SPEED_GRADE     (8),
		.DEV_PACKAGE     (3)
	) axi_adrv9001 (
		.s_axi_aclk                  (sys_hps_h2f_user1_clock_clk),                  //   s_axi_clock.clk
		.s_axi_aresetn               (~rst_controller_reset_out_reset),              //   s_axi_reset.reset_n
		.s_axi_awvalid               (mm_interconnect_0_axi_adrv9001_s_axi_awvalid), //         s_axi.awvalid
		.s_axi_awaddr                (mm_interconnect_0_axi_adrv9001_s_axi_awaddr),  //              .awaddr
		.s_axi_awprot                (mm_interconnect_0_axi_adrv9001_s_axi_awprot),  //              .awprot
		.s_axi_awready               (mm_interconnect_0_axi_adrv9001_s_axi_awready), //              .awready
		.s_axi_wvalid                (mm_interconnect_0_axi_adrv9001_s_axi_wvalid),  //              .wvalid
		.s_axi_wdata                 (mm_interconnect_0_axi_adrv9001_s_axi_wdata),   //              .wdata
		.s_axi_wstrb                 (mm_interconnect_0_axi_adrv9001_s_axi_wstrb),   //              .wstrb
		.s_axi_wready                (mm_interconnect_0_axi_adrv9001_s_axi_wready),  //              .wready
		.s_axi_bvalid                (mm_interconnect_0_axi_adrv9001_s_axi_bvalid),  //              .bvalid
		.s_axi_bresp                 (mm_interconnect_0_axi_adrv9001_s_axi_bresp),   //              .bresp
		.s_axi_bready                (mm_interconnect_0_axi_adrv9001_s_axi_bready),  //              .bready
		.s_axi_arvalid               (mm_interconnect_0_axi_adrv9001_s_axi_arvalid), //              .arvalid
		.s_axi_araddr                (mm_interconnect_0_axi_adrv9001_s_axi_araddr),  //              .araddr
		.s_axi_arprot                (mm_interconnect_0_axi_adrv9001_s_axi_arprot),  //              .arprot
		.s_axi_arready               (mm_interconnect_0_axi_adrv9001_s_axi_arready), //              .arready
		.s_axi_rvalid                (mm_interconnect_0_axi_adrv9001_s_axi_rvalid),  //              .rvalid
		.s_axi_rresp                 (mm_interconnect_0_axi_adrv9001_s_axi_rresp),   //              .rresp
		.s_axi_rdata                 (mm_interconnect_0_axi_adrv9001_s_axi_rdata),   //              .rdata
		.s_axi_rready                (mm_interconnect_0_axi_adrv9001_s_axi_rready),  //              .rready
		.adc_1_clk                   (axi_adrv9001_if_adc_1_clk_clk),                //  if_adc_1_clk.clk
		.adc_2_clk                   (),                                             //  if_adc_2_clk.clk
		.dac_1_clk                   (axi_adrv9001_if_dac_1_clk_clk),                //  if_dac_1_clk.clk
		.dac_2_clk                   (),                                             //  if_dac_2_clk.clk
		.adc_1_rst                   (axi_adrv9001_if_adc_1_rst_reset),              //  if_adc_1_rst.reset
		.adc_2_rst                   (),                                             //  if_adc_2_rst.reset
		.dac_1_rst                   (axi_adrv9001_if_dac_1_rst_reset),              //  if_dac_1_rst.reset
		.dac_2_rst                   (),                                             //  if_dac_2_rst.reset
		.adc_1_enable_i0             (axi_adrv9001_adc_1_ch_0_enable),               //    adc_1_ch_0.enable
		.adc_1_valid_i0              (axi_adrv9001_adc_1_ch_0_valid),                //              .valid
		.adc_1_data_i0               (axi_adrv9001_adc_1_ch_0_data),                 //              .data
		.adc_1_enable_q0             (axi_adrv9001_adc_1_ch_1_enable),               //    adc_1_ch_1.enable
		.adc_1_valid_q0              (axi_adrv9001_adc_1_ch_1_valid),                //              .valid
		.adc_1_data_q0               (axi_adrv9001_adc_1_ch_1_data),                 //              .data
		.adc_1_enable_i1             (axi_adrv9001_adc_1_ch_2_enable),               //    adc_1_ch_2.enable
		.adc_1_valid_i1              (axi_adrv9001_adc_1_ch_2_valid),                //              .valid
		.adc_1_data_i1               (axi_adrv9001_adc_1_ch_2_data),                 //              .data
		.adc_1_enable_q1             (axi_adrv9001_adc_1_ch_3_enable),               //    adc_1_ch_3.enable
		.adc_1_valid_q1              (axi_adrv9001_adc_1_ch_3_valid),                //              .valid
		.adc_1_data_q1               (axi_adrv9001_adc_1_ch_3_data),                 //              .data
		.adc_1_dovf                  (util_adc_wfifo_if_din_ovf_ovf),                // if_adc_1_dovf.ovf
		.adc_2_enable_i0             (),                                             //    adc_2_ch_0.enable
		.adc_2_valid_i0              (),                                             //              .valid
		.adc_2_data_i0               (),                                             //              .data
		.adc_2_enable_q0             (),                                             //    adc_2_ch_1.enable
		.adc_2_valid_q0              (),                                             //              .valid
		.adc_2_data_q0               (),                                             //              .data
		.adc_2_dovf                  (),                                             // if_adc_2_dovf.ovf
		.dac_1_enable_i0             (axi_adrv9001_dac_1_ch_0_enable),               //    dac_1_ch_0.enable
		.dac_1_valid_i0              (axi_adrv9001_dac_1_ch_0_valid),                //              .valid
		.dac_1_data_i0               (util_dac_rfifo_dout_0_data),                   //              .data
		.dac_1_enable_q0             (axi_adrv9001_dac_1_ch_1_enable),               //    dac_1_ch_1.enable
		.dac_1_valid_q0              (axi_adrv9001_dac_1_ch_1_valid),                //              .valid
		.dac_1_data_q0               (util_dac_rfifo_dout_1_data),                   //              .data
		.dac_1_enable_i1             (axi_adrv9001_dac_1_ch_2_enable),               //    dac_1_ch_2.enable
		.dac_1_valid_i1              (axi_adrv9001_dac_1_ch_2_valid),                //              .valid
		.dac_1_data_i1               (util_dac_rfifo_dout_2_data),                   //              .data
		.dac_1_enable_q1             (axi_adrv9001_dac_1_ch_3_enable),               //    dac_1_ch_3.enable
		.dac_1_valid_q1              (axi_adrv9001_dac_1_ch_3_valid),                //              .valid
		.dac_1_data_q1               (util_dac_rfifo_dout_3_data),                   //              .data
		.dac_1_dunf                  (util_dac_rfifo_if_dout_unf_unf),               // if_dac_1_dunf.unf
		.dac_2_enable_i0             (),                                             //    dac_2_ch_0.enable
		.dac_2_valid_i0              (),                                             //              .valid
		.dac_2_data_i0               (),                                             //              .data
		.dac_2_enable_q0             (),                                             //    dac_2_ch_1.enable
		.dac_2_valid_q0              (),                                             //              .valid
		.dac_2_data_q0               (),                                             //              .data
		.dac_2_dunf                  (),                                             // if_dac_2_dunf.unf
		.gpio_rx1_enable_in          (adrv9001_tdd_if_rx1_enable_in),                //        tdd_if.rx1_enable_in
		.gpio_rx2_enable_in          (adrv9001_tdd_if_rx2_enable_in),                //              .rx2_enable_in
		.gpio_tx1_enable_in          (adrv9001_tdd_if_tx1_enable_in),                //              .tx1_enable_in
		.gpio_tx2_enable_in          (adrv9001_tdd_if_tx2_enable_in),                //              .tx2_enable_in
		.tdd_sync                    (adrv9001_tdd_if_tdd_sync_in),                  //              .tdd_sync_in
		.rx1_dclk_in_p_dclk_in       (adrv9001_if_rx1_dclk_in_p_dclk_in),            //     device_if.rx1_dclk_in_p_dclk_in
		.rx1_idata_in_n_idata0       (adrv9001_if_rx1_idata_in_n_idata0),            //              .rx1_idata_in_n_idata0
		.rx1_idata_in_p_idata1       (adrv9001_if_rx1_idata_in_p_idata1),            //              .rx1_idata_in_p_idata1
		.rx1_qdata_in_n_qdata2       (adrv9001_if_rx1_qdata_in_n_qdata2),            //              .rx1_qdata_in_n_qdata2
		.rx1_qdata_in_p_qdata3       (adrv9001_if_rx1_qdata_in_p_qdata3),            //              .rx1_qdata_in_p_qdata3
		.rx1_strobe_in_p_strobe_in   (adrv9001_if_rx1_strobe_in_p_strobe_in),        //              .rx1_strobe_in_p_strobe_in
		.rx1_enable                  (adrv9001_if_rx1_enable),                       //              .rx1_enable
		.rx2_dclk_in_p_dclk_in       (adrv9001_if_rx2_dclk_in_p_dclk_in),            //              .rx2_dclk_in_p_dclk_in
		.rx2_idata_in_n_idata0       (adrv9001_if_rx2_idata_in_n_idata0),            //              .rx2_idata_in_n_idata0
		.rx2_idata_in_p_idata1       (adrv9001_if_rx2_idata_in_p_idata1),            //              .rx2_idata_in_p_idata1
		.rx2_qdata_in_n_qdata2       (adrv9001_if_rx2_qdata_in_n_qdata2),            //              .rx2_qdata_in_n_qdata2
		.rx2_qdata_in_p_qdata3       (adrv9001_if_rx2_qdata_in_p_qdata3),            //              .rx2_qdata_in_p_qdata3
		.rx2_strobe_in_p_strobe_in   (adrv9001_if_rx2_strobe_in_p_strobe_in),        //              .rx2_strobe_in_p_strobe_in
		.rx2_enable                  (adrv9001_if_rx2_enable),                       //              .rx2_enable
		.tx1_dclk_out_p_dclk_out     (adrv9001_if_tx1_dclk_out_p_dclk_out),          //              .tx1_dclk_out_p_dclk_out
		.tx1_dclk_in_p_dclk_in       (adrv9001_if_tx1_dclk_in_p_dclk_in),            //              .tx1_dclk_in_p_dclk_in
		.tx1_idata_out_n_idata0      (adrv9001_if_tx1_idata_out_n_idata0),           //              .tx1_idata_out_n_idata0
		.tx1_idata_out_p_idata1      (adrv9001_if_tx1_idata_out_p_idata1),           //              .tx1_idata_out_p_idata1
		.tx1_qdata_out_n_qdata2      (adrv9001_if_tx1_qdata_out_n_qdata2),           //              .tx1_qdata_out_n_qdata2
		.tx1_qdata_out_p_qdata3      (adrv9001_if_tx1_qdata_out_p_qdata3),           //              .tx1_qdata_out_p_qdata3
		.tx1_strobe_out_p_strobe_out (adrv9001_if_tx1_strobe_out_p_strobe_out),      //              .tx1_strobe_out_p_strobe_out
		.tx1_enable                  (adrv9001_if_tx1_enable),                       //              .tx1_enable
		.tx2_dclk_out_p_dclk_out     (adrv9001_if_tx2_dclk_out_p_dclk_out),          //              .tx2_dclk_out_p_dclk_out
		.tx2_dclk_in_p_dclk_in       (adrv9001_if_tx2_dclk_in_p_dclk_in),            //              .tx2_dclk_in_p_dclk_in
		.tx2_idata_out_n_idata0      (adrv9001_if_tx2_idata_out_n_idata0),           //              .tx2_idata_out_n_idata0
		.tx2_idata_out_p_idata1      (adrv9001_if_tx2_idata_out_p_idata1),           //              .tx2_idata_out_p_idata1
		.tx2_qdata_out_n_qdata2      (adrv9001_if_tx2_qdata_out_n_qdata2),           //              .tx2_qdata_out_n_qdata2
		.tx2_qdata_out_p_qdata3      (adrv9001_if_tx2_qdata_out_p_qdata3),           //              .tx2_qdata_out_p_qdata3
		.tx2_strobe_out_p_strobe_out (adrv9001_if_tx2_strobe_out_p_strobe_out),      //              .tx2_strobe_out_p_strobe_out
		.tx2_enable                  (adrv9001_if_tx2_enable)                        //              .tx2_enable
	);

	axi_dmac #(
		.ID                    (0),
		.DMA_LENGTH_WIDTH      (24),
		.FIFO_SIZE             (4),
		.MAX_BYTES_PER_BURST   (128),
		.DMA_TYPE_SRC          (0),
		.DMA_AXI_PROTOCOL_SRC  (1),
		.DMA_DATA_WIDTH_SRC    (64),
		.AXI_SLICE_SRC         (0),
		.DMA_TYPE_DEST         (1),
		.DMA_AXI_PROTOCOL_DEST (1),
		.DMA_DATA_WIDTH_DEST   (64),
		.AXI_SLICE_DEST        (0),
		.CYCLIC                (1),
		.DMA_2D_TRANSFER       (0),
		.SYNC_TRANSFER_START   (0),
		.ASYNC_CLK_REQ_SRC     (0),
		.ASYNC_CLK_SRC_DEST    (0),
		.ASYNC_CLK_DEST_REQ    (0),
		.ENABLE_DIAGNOSTICS_IF (0),
		.DMA_AXIS_ID_W         (8),
		.DMA_AXIS_DEST_W       (4)
	) axi_dac_dma (
		.s_axi_aclk             (sys_hps_h2f_user1_clock_clk),                                          //        s_axi_clock.clk
		.s_axi_aresetn          (~rst_controller_reset_out_reset),                                      //        s_axi_reset.reset_n
		.s_axi_awvalid          (mm_interconnect_0_axi_dac_dma_s_axi_awvalid),                          //              s_axi.awvalid
		.s_axi_awaddr           (mm_interconnect_0_axi_dac_dma_s_axi_awaddr),                           //                   .awaddr
		.s_axi_awprot           (mm_interconnect_0_axi_dac_dma_s_axi_awprot),                           //                   .awprot
		.s_axi_awready          (mm_interconnect_0_axi_dac_dma_s_axi_awready),                          //                   .awready
		.s_axi_wvalid           (mm_interconnect_0_axi_dac_dma_s_axi_wvalid),                           //                   .wvalid
		.s_axi_wdata            (mm_interconnect_0_axi_dac_dma_s_axi_wdata),                            //                   .wdata
		.s_axi_wstrb            (mm_interconnect_0_axi_dac_dma_s_axi_wstrb),                            //                   .wstrb
		.s_axi_wready           (mm_interconnect_0_axi_dac_dma_s_axi_wready),                           //                   .wready
		.s_axi_bvalid           (mm_interconnect_0_axi_dac_dma_s_axi_bvalid),                           //                   .bvalid
		.s_axi_bresp            (mm_interconnect_0_axi_dac_dma_s_axi_bresp),                            //                   .bresp
		.s_axi_bready           (mm_interconnect_0_axi_dac_dma_s_axi_bready),                           //                   .bready
		.s_axi_arvalid          (mm_interconnect_0_axi_dac_dma_s_axi_arvalid),                          //                   .arvalid
		.s_axi_araddr           (mm_interconnect_0_axi_dac_dma_s_axi_araddr),                           //                   .araddr
		.s_axi_arprot           (mm_interconnect_0_axi_dac_dma_s_axi_arprot),                           //                   .arprot
		.s_axi_arready          (mm_interconnect_0_axi_dac_dma_s_axi_arready),                          //                   .arready
		.s_axi_rvalid           (mm_interconnect_0_axi_dac_dma_s_axi_rvalid),                           //                   .rvalid
		.s_axi_rresp            (mm_interconnect_0_axi_dac_dma_s_axi_rresp),                            //                   .rresp
		.s_axi_rdata            (mm_interconnect_0_axi_dac_dma_s_axi_rdata),                            //                   .rdata
		.s_axi_rready           (mm_interconnect_0_axi_dac_dma_s_axi_rready),                           //                   .rready
		.irq                    (irq_mapper_receiver2_irq),                                             //   interrupt_sender.irq
		.m_src_axi_aclk         (sys_hps_h2f_user1_clock_clk),                                          //    m_src_axi_clock.clk
		.m_src_axi_aresetn      (~rst_controller_reset_out_reset),                                      //    m_src_axi_reset.reset_n
		.m_axis_aclk            (sys_hps_h2f_user1_clock_clk),                                          //     if_m_axis_aclk.clk
		.m_axis_xfer_req        (),                                                                     // if_m_axis_xfer_req.xfer_req
		.m_axis_valid           (axi_dac_dma_m_axis_tvalid),                                            //             m_axis.tvalid
		.m_axis_ready           (axi_dac_dma_m_axis_tready),                                            //                   .tready
		.m_axis_data            (axi_dac_dma_m_axis_tdata),                                             //                   .tdata
		.m_src_axi_awvalid      (axi_dac_dma_m_src_axi_awvalid),                                        //          m_src_axi.awvalid
		.m_src_axi_awaddr       (axi_dac_dma_m_src_axi_awaddr),                                         //                   .awaddr
		.m_src_axi_awready      (axi_dac_dma_m_src_axi_awready),                                        //                   .awready
		.m_src_axi_wvalid       (axi_dac_dma_m_src_axi_wvalid),                                         //                   .wvalid
		.m_src_axi_wdata        (axi_dac_dma_m_src_axi_wdata),                                          //                   .wdata
		.m_src_axi_wstrb        (axi_dac_dma_m_src_axi_wstrb),                                          //                   .wstrb
		.m_src_axi_wready       (axi_dac_dma_m_src_axi_wready),                                         //                   .wready
		.m_src_axi_bvalid       (axi_dac_dma_m_src_axi_bvalid),                                         //                   .bvalid
		.m_src_axi_bresp        (axi_dac_dma_m_src_axi_bresp),                                          //                   .bresp
		.m_src_axi_bready       (axi_dac_dma_m_src_axi_bready),                                         //                   .bready
		.m_src_axi_arvalid      (axi_dac_dma_m_src_axi_arvalid),                                        //                   .arvalid
		.m_src_axi_araddr       (axi_dac_dma_m_src_axi_araddr),                                         //                   .araddr
		.m_src_axi_arready      (axi_dac_dma_m_src_axi_arready),                                        //                   .arready
		.m_src_axi_rvalid       (axi_dac_dma_m_src_axi_rvalid),                                         //                   .rvalid
		.m_src_axi_rresp        (axi_dac_dma_m_src_axi_rresp),                                          //                   .rresp
		.m_src_axi_rdata        (axi_dac_dma_m_src_axi_rdata),                                          //                   .rdata
		.m_src_axi_rready       (axi_dac_dma_m_src_axi_rready),                                         //                   .rready
		.m_src_axi_awlen        (axi_dac_dma_m_src_axi_awlen),                                          //                   .awlen
		.m_src_axi_awsize       (axi_dac_dma_m_src_axi_awsize),                                         //                   .awsize
		.m_src_axi_awburst      (axi_dac_dma_m_src_axi_awburst),                                        //                   .awburst
		.m_src_axi_awcache      (axi_dac_dma_m_src_axi_awcache),                                        //                   .awcache
		.m_src_axi_awprot       (axi_dac_dma_m_src_axi_awprot),                                         //                   .awprot
		.m_src_axi_wlast        (axi_dac_dma_m_src_axi_wlast),                                          //                   .wlast
		.m_src_axi_arlen        (axi_dac_dma_m_src_axi_arlen),                                          //                   .arlen
		.m_src_axi_arsize       (axi_dac_dma_m_src_axi_arsize),                                         //                   .arsize
		.m_src_axi_arburst      (axi_dac_dma_m_src_axi_arburst),                                        //                   .arburst
		.m_src_axi_arcache      (axi_dac_dma_m_src_axi_arcache),                                        //                   .arcache
		.m_src_axi_arprot       (axi_dac_dma_m_src_axi_arprot),                                         //                   .arprot
		.m_src_axi_awid         (axi_dac_dma_m_src_axi_awid),                                           //                   .awid
		.m_src_axi_awlock       (axi_dac_dma_m_src_axi_awlock),                                         //                   .awlock
		.m_src_axi_wid          (axi_dac_dma_m_src_axi_wid),                                            //                   .wid
		.m_src_axi_arid         (axi_dac_dma_m_src_axi_arid),                                           //                   .arid
		.m_src_axi_arlock       (axi_dac_dma_m_src_axi_arlock),                                         //                   .arlock
		.m_src_axi_rid          (axi_dac_dma_m_src_axi_rid),                                            //                   .rid
		.m_src_axi_bid          (axi_dac_dma_m_src_axi_bid),                                            //                   .bid
		.m_src_axi_rlast        (axi_dac_dma_m_src_axi_rlast),                                          //                   .rlast
		.m_axis_last            (),                                                                     //        (terminated)
		.m_axis_user            (),                                                                     //        (terminated)
		.m_axis_id              (),                                                                     //        (terminated)
		.m_axis_dest            (),                                                                     //        (terminated)
		.m_axis_strb            (),                                                                     //        (terminated)
		.m_axis_keep            (),                                                                     //        (terminated)
		.m_dest_axi_aclk        (1'b0),                                                                 //        (terminated)
		.m_dest_axi_aresetn     (1'b1),                                                                 //        (terminated)
		.s_axis_aclk            (1'b0),                                                                 //        (terminated)
		.s_axis_xfer_req        (),                                                                     //        (terminated)
		.s_axis_valid           (1'b0),                                                                 //        (terminated)
		.s_axis_last            (1'b0),                                                                 //        (terminated)
		.s_axis_ready           (),                                                                     //        (terminated)
		.s_axis_data            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.s_axis_user            (1'b0),                                                                 //        (terminated)
		.s_axis_id              (8'b00000000),                                                          //        (terminated)
		.s_axis_dest            (4'b0000),                                                              //        (terminated)
		.s_axis_strb            (8'b00000000),                                                          //        (terminated)
		.s_axis_keep            (8'b00000000),                                                          //        (terminated)
		.fifo_rd_clk            (1'b0),                                                                 //        (terminated)
		.fifo_rd_en             (1'b0),                                                                 //        (terminated)
		.fifo_rd_valid          (),                                                                     //        (terminated)
		.fifo_rd_dout           (),                                                                     //        (terminated)
		.fifo_rd_underflow      (),                                                                     //        (terminated)
		.fifo_rd_xfer_req       (),                                                                     //        (terminated)
		.fifo_wr_clk            (1'b0),                                                                 //        (terminated)
		.fifo_wr_en             (1'b0),                                                                 //        (terminated)
		.fifo_wr_din            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.fifo_wr_overflow       (),                                                                     //        (terminated)
		.fifo_wr_sync           (1'b0),                                                                 //        (terminated)
		.fifo_wr_xfer_req       (),                                                                     //        (terminated)
		.dest_diag_level_bursts (),                                                                     //        (terminated)
		.m_dest_axi_awvalid     (),                                                                     //        (terminated)
		.m_dest_axi_awaddr      (),                                                                     //        (terminated)
		.m_dest_axi_awready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_wvalid      (),                                                                     //        (terminated)
		.m_dest_axi_wdata       (),                                                                     //        (terminated)
		.m_dest_axi_wstrb       (),                                                                     //        (terminated)
		.m_dest_axi_wready      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_bready      (),                                                                     //        (terminated)
		.m_dest_axi_arvalid     (),                                                                     //        (terminated)
		.m_dest_axi_araddr      (),                                                                     //        (terminated)
		.m_dest_axi_arready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_rdata       (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.m_dest_axi_rready      (),                                                                     //        (terminated)
		.m_dest_axi_awlen       (),                                                                     //        (terminated)
		.m_dest_axi_awsize      (),                                                                     //        (terminated)
		.m_dest_axi_awburst     (),                                                                     //        (terminated)
		.m_dest_axi_awcache     (),                                                                     //        (terminated)
		.m_dest_axi_awprot      (),                                                                     //        (terminated)
		.m_dest_axi_wlast       (),                                                                     //        (terminated)
		.m_dest_axi_arlen       (),                                                                     //        (terminated)
		.m_dest_axi_arsize      (),                                                                     //        (terminated)
		.m_dest_axi_arburst     (),                                                                     //        (terminated)
		.m_dest_axi_arcache     (),                                                                     //        (terminated)
		.m_dest_axi_arprot      (),                                                                     //        (terminated)
		.m_dest_axi_awid        (),                                                                     //        (terminated)
		.m_dest_axi_awlock      (),                                                                     //        (terminated)
		.m_dest_axi_wid         (),                                                                     //        (terminated)
		.m_dest_axi_arid        (),                                                                     //        (terminated)
		.m_dest_axi_arlock      (),                                                                     //        (terminated)
		.m_dest_axi_rid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rlast       (1'b0)                                                                  //        (terminated)
	);

	axi_hdmi_tx #(
		.ID               (0),
		.FPGA_TECHNOLOGY  (101),
		.INTERFACE        ("16_BIT"),
		.CR_CB_N          (0),
		.OUT_CLK_POLARITY (0)
	) axi_hdmi_tx_0 (
		.s_axi_aclk        (sys_hps_h2f_user1_clock_clk),                   // s_axi_clock.clk
		.s_axi_awvalid     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awvalid), //       s_axi.awvalid
		.s_axi_awaddr      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awaddr),  //            .awaddr
		.s_axi_awprot      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awprot),  //            .awprot
		.s_axi_awready     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awready), //            .awready
		.s_axi_wvalid      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wvalid),  //            .wvalid
		.s_axi_wdata       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wdata),   //            .wdata
		.s_axi_wstrb       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wstrb),   //            .wstrb
		.s_axi_wready      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wready),  //            .wready
		.s_axi_bvalid      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bvalid),  //            .bvalid
		.s_axi_bresp       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bresp),   //            .bresp
		.s_axi_bready      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bready),  //            .bready
		.s_axi_arvalid     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arvalid), //            .arvalid
		.s_axi_araddr      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_araddr),  //            .araddr
		.s_axi_arprot      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arprot),  //            .arprot
		.s_axi_arready     (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arready), //            .arready
		.s_axi_rvalid      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rvalid),  //            .rvalid
		.s_axi_rresp       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rresp),   //            .rresp
		.s_axi_rdata       (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rdata),   //            .rdata
		.s_axi_rready      (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rready),  //            .rready
		.hdmi_clk          (hdmi_pll_outclk0_clk),                          //  hdmi_clock.clk
		.hdmi_out_clk      (hdmi_out_h_clk),                                //     hdmi_if.h_clk
		.hdmi_16_hsync     (hdmi_out_h16_hsync),                            //            .h16_hsync
		.hdmi_16_vsync     (hdmi_out_h16_vsync),                            //            .h16_vsync
		.hdmi_16_data_e    (hdmi_out_h16_data_e),                           //            .h16_data_e
		.hdmi_16_data      (hdmi_out_h16_data),                             //            .h16_data
		.hdmi_16_es_data   (hdmi_out_h16_es_data),                          //            .h16_es_data
		.hdmi_24_hsync     (hdmi_out_h24_hsync),                            //            .h24_hsync
		.hdmi_24_vsync     (hdmi_out_h24_vsync),                            //            .h24_vsync
		.hdmi_24_data_e    (hdmi_out_h24_data_e),                           //            .h24_data_e
		.hdmi_24_data      (hdmi_out_h24_data),                             //            .h24_data
		.hdmi_36_hsync     (hdmi_out_h36_hsync),                            //            .h36_hsync
		.hdmi_36_vsync     (hdmi_out_h36_vsync),                            //            .h36_vsync
		.hdmi_36_data_e    (hdmi_out_h36_data_e),                           //            .h36_data_e
		.hdmi_36_data      (hdmi_out_h36_data),                             //            .h36_data
		.vdma_clk          (sys_hps_h2f_user1_clock_clk),                   //  vdma_clock.clk
		.s_axi_aresetn     (~rst_controller_reset_out_reset),               //  vdma_reset.reset_n
		.vdma_end_of_frame (hdmi_dmac_0_m_axis_tlast),                      //     vdma_if.tlast
		.vdma_valid        (hdmi_dmac_0_m_axis_tvalid),                     //            .tvalid
		.vdma_data         (hdmi_dmac_0_m_axis_tdata),                      //            .tdata
		.vdma_ready        (hdmi_dmac_0_m_axis_tready)                      //            .tready
	);

	axi_dmac #(
		.ID                    (0),
		.DMA_LENGTH_WIDTH      (24),
		.FIFO_SIZE             (8),
		.MAX_BYTES_PER_BURST   (128),
		.DMA_TYPE_SRC          (0),
		.DMA_AXI_PROTOCOL_SRC  (1),
		.DMA_DATA_WIDTH_SRC    (64),
		.AXI_SLICE_SRC         (0),
		.DMA_TYPE_DEST         (1),
		.DMA_AXI_PROTOCOL_DEST (1),
		.DMA_DATA_WIDTH_DEST   (64),
		.AXI_SLICE_DEST        (0),
		.CYCLIC                (1),
		.DMA_2D_TRANSFER       (1),
		.SYNC_TRANSFER_START   (0),
		.ASYNC_CLK_REQ_SRC     (0),
		.ASYNC_CLK_SRC_DEST    (0),
		.ASYNC_CLK_DEST_REQ    (0),
		.ENABLE_DIAGNOSTICS_IF (0),
		.DMA_AXIS_ID_W         (8),
		.DMA_AXIS_DEST_W       (4)
	) hdmi_dmac_0 (
		.s_axi_aclk             (sys_hps_h2f_user1_clock_clk),                                          //        s_axi_clock.clk
		.s_axi_aresetn          (~rst_controller_reset_out_reset),                                      //        s_axi_reset.reset_n
		.s_axi_awvalid          (mm_interconnect_0_hdmi_dmac_0_s_axi_awvalid),                          //              s_axi.awvalid
		.s_axi_awaddr           (mm_interconnect_0_hdmi_dmac_0_s_axi_awaddr),                           //                   .awaddr
		.s_axi_awprot           (mm_interconnect_0_hdmi_dmac_0_s_axi_awprot),                           //                   .awprot
		.s_axi_awready          (mm_interconnect_0_hdmi_dmac_0_s_axi_awready),                          //                   .awready
		.s_axi_wvalid           (mm_interconnect_0_hdmi_dmac_0_s_axi_wvalid),                           //                   .wvalid
		.s_axi_wdata            (mm_interconnect_0_hdmi_dmac_0_s_axi_wdata),                            //                   .wdata
		.s_axi_wstrb            (mm_interconnect_0_hdmi_dmac_0_s_axi_wstrb),                            //                   .wstrb
		.s_axi_wready           (mm_interconnect_0_hdmi_dmac_0_s_axi_wready),                           //                   .wready
		.s_axi_bvalid           (mm_interconnect_0_hdmi_dmac_0_s_axi_bvalid),                           //                   .bvalid
		.s_axi_bresp            (mm_interconnect_0_hdmi_dmac_0_s_axi_bresp),                            //                   .bresp
		.s_axi_bready           (mm_interconnect_0_hdmi_dmac_0_s_axi_bready),                           //                   .bready
		.s_axi_arvalid          (mm_interconnect_0_hdmi_dmac_0_s_axi_arvalid),                          //                   .arvalid
		.s_axi_araddr           (mm_interconnect_0_hdmi_dmac_0_s_axi_araddr),                           //                   .araddr
		.s_axi_arprot           (mm_interconnect_0_hdmi_dmac_0_s_axi_arprot),                           //                   .arprot
		.s_axi_arready          (mm_interconnect_0_hdmi_dmac_0_s_axi_arready),                          //                   .arready
		.s_axi_rvalid           (mm_interconnect_0_hdmi_dmac_0_s_axi_rvalid),                           //                   .rvalid
		.s_axi_rresp            (mm_interconnect_0_hdmi_dmac_0_s_axi_rresp),                            //                   .rresp
		.s_axi_rdata            (mm_interconnect_0_hdmi_dmac_0_s_axi_rdata),                            //                   .rdata
		.s_axi_rready           (mm_interconnect_0_hdmi_dmac_0_s_axi_rready),                           //                   .rready
		.irq                    (irq_mapper_receiver0_irq),                                             //   interrupt_sender.irq
		.m_src_axi_aclk         (sys_hps_h2f_user1_clock_clk),                                          //    m_src_axi_clock.clk
		.m_src_axi_aresetn      (~rst_controller_reset_out_reset),                                      //    m_src_axi_reset.reset_n
		.m_axis_aclk            (sys_hps_h2f_user1_clock_clk),                                          //     if_m_axis_aclk.clk
		.m_axis_xfer_req        (),                                                                     // if_m_axis_xfer_req.xfer_req
		.m_axis_valid           (hdmi_dmac_0_m_axis_tvalid),                                            //             m_axis.tvalid
		.m_axis_last            (hdmi_dmac_0_m_axis_tlast),                                             //                   .tlast
		.m_axis_ready           (hdmi_dmac_0_m_axis_tready),                                            //                   .tready
		.m_axis_data            (hdmi_dmac_0_m_axis_tdata),                                             //                   .tdata
		.m_src_axi_awvalid      (hdmi_dmac_0_m_src_axi_awvalid),                                        //          m_src_axi.awvalid
		.m_src_axi_awaddr       (hdmi_dmac_0_m_src_axi_awaddr),                                         //                   .awaddr
		.m_src_axi_awready      (hdmi_dmac_0_m_src_axi_awready),                                        //                   .awready
		.m_src_axi_wvalid       (hdmi_dmac_0_m_src_axi_wvalid),                                         //                   .wvalid
		.m_src_axi_wdata        (hdmi_dmac_0_m_src_axi_wdata),                                          //                   .wdata
		.m_src_axi_wstrb        (hdmi_dmac_0_m_src_axi_wstrb),                                          //                   .wstrb
		.m_src_axi_wready       (hdmi_dmac_0_m_src_axi_wready),                                         //                   .wready
		.m_src_axi_bvalid       (hdmi_dmac_0_m_src_axi_bvalid),                                         //                   .bvalid
		.m_src_axi_bresp        (hdmi_dmac_0_m_src_axi_bresp),                                          //                   .bresp
		.m_src_axi_bready       (hdmi_dmac_0_m_src_axi_bready),                                         //                   .bready
		.m_src_axi_arvalid      (hdmi_dmac_0_m_src_axi_arvalid),                                        //                   .arvalid
		.m_src_axi_araddr       (hdmi_dmac_0_m_src_axi_araddr),                                         //                   .araddr
		.m_src_axi_arready      (hdmi_dmac_0_m_src_axi_arready),                                        //                   .arready
		.m_src_axi_rvalid       (hdmi_dmac_0_m_src_axi_rvalid),                                         //                   .rvalid
		.m_src_axi_rresp        (hdmi_dmac_0_m_src_axi_rresp),                                          //                   .rresp
		.m_src_axi_rdata        (hdmi_dmac_0_m_src_axi_rdata),                                          //                   .rdata
		.m_src_axi_rready       (hdmi_dmac_0_m_src_axi_rready),                                         //                   .rready
		.m_src_axi_awlen        (hdmi_dmac_0_m_src_axi_awlen),                                          //                   .awlen
		.m_src_axi_awsize       (hdmi_dmac_0_m_src_axi_awsize),                                         //                   .awsize
		.m_src_axi_awburst      (hdmi_dmac_0_m_src_axi_awburst),                                        //                   .awburst
		.m_src_axi_awcache      (hdmi_dmac_0_m_src_axi_awcache),                                        //                   .awcache
		.m_src_axi_awprot       (hdmi_dmac_0_m_src_axi_awprot),                                         //                   .awprot
		.m_src_axi_wlast        (hdmi_dmac_0_m_src_axi_wlast),                                          //                   .wlast
		.m_src_axi_arlen        (hdmi_dmac_0_m_src_axi_arlen),                                          //                   .arlen
		.m_src_axi_arsize       (hdmi_dmac_0_m_src_axi_arsize),                                         //                   .arsize
		.m_src_axi_arburst      (hdmi_dmac_0_m_src_axi_arburst),                                        //                   .arburst
		.m_src_axi_arcache      (hdmi_dmac_0_m_src_axi_arcache),                                        //                   .arcache
		.m_src_axi_arprot       (hdmi_dmac_0_m_src_axi_arprot),                                         //                   .arprot
		.m_src_axi_awid         (hdmi_dmac_0_m_src_axi_awid),                                           //                   .awid
		.m_src_axi_awlock       (hdmi_dmac_0_m_src_axi_awlock),                                         //                   .awlock
		.m_src_axi_wid          (hdmi_dmac_0_m_src_axi_wid),                                            //                   .wid
		.m_src_axi_arid         (hdmi_dmac_0_m_src_axi_arid),                                           //                   .arid
		.m_src_axi_arlock       (hdmi_dmac_0_m_src_axi_arlock),                                         //                   .arlock
		.m_src_axi_rid          (hdmi_dmac_0_m_src_axi_rid),                                            //                   .rid
		.m_src_axi_bid          (hdmi_dmac_0_m_src_axi_bid),                                            //                   .bid
		.m_src_axi_rlast        (hdmi_dmac_0_m_src_axi_rlast),                                          //                   .rlast
		.m_axis_user            (),                                                                     //        (terminated)
		.m_axis_id              (),                                                                     //        (terminated)
		.m_axis_dest            (),                                                                     //        (terminated)
		.m_axis_strb            (),                                                                     //        (terminated)
		.m_axis_keep            (),                                                                     //        (terminated)
		.m_dest_axi_aclk        (1'b0),                                                                 //        (terminated)
		.m_dest_axi_aresetn     (1'b1),                                                                 //        (terminated)
		.s_axis_aclk            (1'b0),                                                                 //        (terminated)
		.s_axis_xfer_req        (),                                                                     //        (terminated)
		.s_axis_valid           (1'b0),                                                                 //        (terminated)
		.s_axis_last            (1'b0),                                                                 //        (terminated)
		.s_axis_ready           (),                                                                     //        (terminated)
		.s_axis_data            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.s_axis_user            (1'b0),                                                                 //        (terminated)
		.s_axis_id              (8'b00000000),                                                          //        (terminated)
		.s_axis_dest            (4'b0000),                                                              //        (terminated)
		.s_axis_strb            (8'b00000000),                                                          //        (terminated)
		.s_axis_keep            (8'b00000000),                                                          //        (terminated)
		.fifo_rd_clk            (1'b0),                                                                 //        (terminated)
		.fifo_rd_en             (1'b0),                                                                 //        (terminated)
		.fifo_rd_valid          (),                                                                     //        (terminated)
		.fifo_rd_dout           (),                                                                     //        (terminated)
		.fifo_rd_underflow      (),                                                                     //        (terminated)
		.fifo_rd_xfer_req       (),                                                                     //        (terminated)
		.fifo_wr_clk            (1'b0),                                                                 //        (terminated)
		.fifo_wr_en             (1'b0),                                                                 //        (terminated)
		.fifo_wr_din            (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.fifo_wr_overflow       (),                                                                     //        (terminated)
		.fifo_wr_sync           (1'b0),                                                                 //        (terminated)
		.fifo_wr_xfer_req       (),                                                                     //        (terminated)
		.dest_diag_level_bursts (),                                                                     //        (terminated)
		.m_dest_axi_awvalid     (),                                                                     //        (terminated)
		.m_dest_axi_awaddr      (),                                                                     //        (terminated)
		.m_dest_axi_awready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_wvalid      (),                                                                     //        (terminated)
		.m_dest_axi_wdata       (),                                                                     //        (terminated)
		.m_dest_axi_wstrb       (),                                                                     //        (terminated)
		.m_dest_axi_wready      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_bready      (),                                                                     //        (terminated)
		.m_dest_axi_arvalid     (),                                                                     //        (terminated)
		.m_dest_axi_araddr      (),                                                                     //        (terminated)
		.m_dest_axi_arready     (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rvalid      (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rresp       (2'b00),                                                                //        (terminated)
		.m_dest_axi_rdata       (64'b0000000000000000000000000000000000000000000000000000000000000000), //        (terminated)
		.m_dest_axi_rready      (),                                                                     //        (terminated)
		.m_dest_axi_awlen       (),                                                                     //        (terminated)
		.m_dest_axi_awsize      (),                                                                     //        (terminated)
		.m_dest_axi_awburst     (),                                                                     //        (terminated)
		.m_dest_axi_awcache     (),                                                                     //        (terminated)
		.m_dest_axi_awprot      (),                                                                     //        (terminated)
		.m_dest_axi_wlast       (),                                                                     //        (terminated)
		.m_dest_axi_arlen       (),                                                                     //        (terminated)
		.m_dest_axi_arsize      (),                                                                     //        (terminated)
		.m_dest_axi_arburst     (),                                                                     //        (terminated)
		.m_dest_axi_arcache     (),                                                                     //        (terminated)
		.m_dest_axi_arprot      (),                                                                     //        (terminated)
		.m_dest_axi_awid        (),                                                                     //        (terminated)
		.m_dest_axi_awlock      (),                                                                     //        (terminated)
		.m_dest_axi_wid         (),                                                                     //        (terminated)
		.m_dest_axi_arid        (),                                                                     //        (terminated)
		.m_dest_axi_arlock      (),                                                                     //        (terminated)
		.m_dest_axi_rid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_bid         (1'b0),                                                                 //        (terminated)
		.m_dest_axi_rlast       (1'b0)                                                                  //        (terminated)
	);

	system_bd_hdmi_pll hdmi_pll (
		.refclk   (sys_hps_h2f_user1_clock_clk), //  refclk.clk
		.rst      (~sys_rst_reset_n),            //   reset.reset
		.outclk_0 (hdmi_pll_outclk0_clk),        // outclk0.clk
		.locked   ()                             // (terminated)
	);

	system_bd_spi_0 spi_0 (
		.clk           (sys_hps_h2f_user1_clock_clk),                         //              clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver5_irq),                            //              irq.irq
		.MISO          (spi_0_external_MISO),                                 //         external.export
		.MOSI          (spi_0_external_MOSI),                                 //                 .export
		.SCLK          (spi_0_external_SCLK),                                 //                 .export
		.SS_n          (spi_0_external_SS_n)                                  //                 .export
	);

	system_bd_sys_gpio_bd sys_gpio_bd (
		.clk        (sys_hps_h2f_user1_clock_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_bd_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_bd_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_bd_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_bd_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_bd_s1_readdata),   //                    .readdata
		.in_port    (sys_gpio_bd_in_port),                         // external_connection.export
		.out_port   (sys_gpio_bd_out_port),                        //                    .export
		.irq        (irq_mapper_receiver3_irq)                     //                 irq.irq
	);

	system_bd_sys_gpio_in sys_gpio_in (
		.clk        (sys_hps_h2f_user1_clock_clk),                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_in_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_in_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_in_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_in_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_in_s1_readdata),   //                    .readdata
		.in_port    (sys_gpio_in_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                     //                 irq.irq
	);

	system_bd_sys_gpio_out sys_gpio_out (
		.clk        (sys_hps_h2f_user1_clock_clk),                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_sys_gpio_out_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sys_gpio_out_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sys_gpio_out_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sys_gpio_out_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sys_gpio_out_s1_readdata),   //                    .readdata
		.out_port   (sys_gpio_out_export)                           // external_connection.export
	);

	system_bd_sys_hps #(
		.F2S_Width (2),
		.S2F_Width (2)
	) sys_hps (
		.h2f_user1_clk            (sys_hps_h2f_user1_clock_clk),                             //   h2f_user1_clock.clk
		.mem_a                    (sys_hps_memory_mem_a),                                    //            memory.mem_a
		.mem_ba                   (sys_hps_memory_mem_ba),                                   //                  .mem_ba
		.mem_ck                   (sys_hps_memory_mem_ck),                                   //                  .mem_ck
		.mem_ck_n                 (sys_hps_memory_mem_ck_n),                                 //                  .mem_ck_n
		.mem_cke                  (sys_hps_memory_mem_cke),                                  //                  .mem_cke
		.mem_cs_n                 (sys_hps_memory_mem_cs_n),                                 //                  .mem_cs_n
		.mem_ras_n                (sys_hps_memory_mem_ras_n),                                //                  .mem_ras_n
		.mem_cas_n                (sys_hps_memory_mem_cas_n),                                //                  .mem_cas_n
		.mem_we_n                 (sys_hps_memory_mem_we_n),                                 //                  .mem_we_n
		.mem_reset_n              (sys_hps_memory_mem_reset_n),                              //                  .mem_reset_n
		.mem_dq                   (sys_hps_memory_mem_dq),                                   //                  .mem_dq
		.mem_dqs                  (sys_hps_memory_mem_dqs),                                  //                  .mem_dqs
		.mem_dqs_n                (sys_hps_memory_mem_dqs_n),                                //                  .mem_dqs_n
		.mem_odt                  (sys_hps_memory_mem_odt),                                  //                  .mem_odt
		.mem_dm                   (sys_hps_memory_mem_dm),                                   //                  .mem_dm
		.oct_rzqin                (sys_hps_memory_oct_rzqin),                                //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (sys_hps_hps_io_hps_io_emac1_inst_TX_CLK),                 //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (sys_hps_hps_io_hps_io_emac1_inst_TXD0),                   //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (sys_hps_hps_io_hps_io_emac1_inst_TXD1),                   //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (sys_hps_hps_io_hps_io_emac1_inst_TXD2),                   //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (sys_hps_hps_io_hps_io_emac1_inst_TXD3),                   //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (sys_hps_hps_io_hps_io_emac1_inst_RXD0),                   //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (sys_hps_hps_io_hps_io_emac1_inst_MDIO),                   //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (sys_hps_hps_io_hps_io_emac1_inst_MDC),                    //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (sys_hps_hps_io_hps_io_emac1_inst_RX_CTL),                 //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (sys_hps_hps_io_hps_io_emac1_inst_TX_CTL),                 //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (sys_hps_hps_io_hps_io_emac1_inst_RX_CLK),                 //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (sys_hps_hps_io_hps_io_emac1_inst_RXD1),                   //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (sys_hps_hps_io_hps_io_emac1_inst_RXD2),                   //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (sys_hps_hps_io_hps_io_emac1_inst_RXD3),                   //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (sys_hps_hps_io_hps_io_qspi_inst_IO0),                     //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (sys_hps_hps_io_hps_io_qspi_inst_IO1),                     //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (sys_hps_hps_io_hps_io_qspi_inst_IO2),                     //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (sys_hps_hps_io_hps_io_qspi_inst_IO3),                     //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (sys_hps_hps_io_hps_io_qspi_inst_SS0),                     //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (sys_hps_hps_io_hps_io_qspi_inst_CLK),                     //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (sys_hps_hps_io_hps_io_sdio_inst_CMD),                     //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (sys_hps_hps_io_hps_io_sdio_inst_D0),                      //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (sys_hps_hps_io_hps_io_sdio_inst_D1),                      //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (sys_hps_hps_io_hps_io_sdio_inst_CLK),                     //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (sys_hps_hps_io_hps_io_sdio_inst_D2),                      //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (sys_hps_hps_io_hps_io_sdio_inst_D3),                      //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (sys_hps_hps_io_hps_io_usb1_inst_D0),                      //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (sys_hps_hps_io_hps_io_usb1_inst_D1),                      //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (sys_hps_hps_io_hps_io_usb1_inst_D2),                      //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (sys_hps_hps_io_hps_io_usb1_inst_D3),                      //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (sys_hps_hps_io_hps_io_usb1_inst_D4),                      //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (sys_hps_hps_io_hps_io_usb1_inst_D5),                      //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (sys_hps_hps_io_hps_io_usb1_inst_D6),                      //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (sys_hps_hps_io_hps_io_usb1_inst_D7),                      //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (sys_hps_hps_io_hps_io_usb1_inst_CLK),                     //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (sys_hps_hps_io_hps_io_usb1_inst_STP),                     //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (sys_hps_hps_io_hps_io_usb1_inst_DIR),                     //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (sys_hps_hps_io_hps_io_usb1_inst_NXT),                     //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (sys_hps_hps_io_hps_io_uart0_inst_RX),                     //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (sys_hps_hps_io_hps_io_uart0_inst_TX),                     //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (sys_hps_hps_io_hps_io_i2c0_inst_SDA),                     //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (sys_hps_hps_io_hps_io_i2c0_inst_SCL),                     //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (sys_hps_hps_io_hps_io_i2c1_inst_SDA),                     //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (sys_hps_hps_io_hps_io_i2c1_inst_SCL),                     //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO00  (sys_hps_hps_io_hps_io_gpio_inst_GPIO00),                  //                  .hps_io_gpio_inst_GPIO00
		.hps_io_gpio_inst_GPIO09  (sys_hps_hps_io_hps_io_gpio_inst_GPIO09),                  //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (sys_hps_hps_io_hps_io_gpio_inst_GPIO35),                  //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (sys_hps_hps_io_hps_io_gpio_inst_GPIO40),                  //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (sys_hps_hps_io_hps_io_gpio_inst_GPIO41),                  //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO42  (sys_hps_hps_io_hps_io_gpio_inst_GPIO42),                  //                  .hps_io_gpio_inst_GPIO42
		.hps_io_gpio_inst_GPIO43  (sys_hps_hps_io_hps_io_gpio_inst_GPIO43),                  //                  .hps_io_gpio_inst_GPIO43
		.hps_io_gpio_inst_GPIO44  (sys_hps_hps_io_hps_io_gpio_inst_GPIO44),                  //                  .hps_io_gpio_inst_GPIO44
		.hps_io_gpio_inst_GPIO48  (sys_hps_hps_io_hps_io_gpio_inst_GPIO48),                  //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (sys_hps_hps_io_hps_io_gpio_inst_GPIO53),                  //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (sys_hps_hps_io_hps_io_gpio_inst_GPIO54),                  //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO55  (sys_hps_hps_io_hps_io_gpio_inst_GPIO55),                  //                  .hps_io_gpio_inst_GPIO55
		.hps_io_gpio_inst_GPIO56  (sys_hps_hps_io_hps_io_gpio_inst_GPIO56),                  //                  .hps_io_gpio_inst_GPIO56
		.hps_io_gpio_inst_GPIO57  (sys_hps_hps_io_hps_io_gpio_inst_GPIO57),                  //                  .hps_io_gpio_inst_GPIO57
		.hps_io_gpio_inst_GPIO58  (sys_hps_hps_io_hps_io_gpio_inst_GPIO58),                  //                  .hps_io_gpio_inst_GPIO58
		.hps_io_gpio_inst_GPIO59  (sys_hps_hps_io_hps_io_gpio_inst_GPIO59),                  //                  .hps_io_gpio_inst_GPIO59
		.hps_io_gpio_inst_GPIO61  (sys_hps_hps_io_hps_io_gpio_inst_GPIO61),                  //                  .hps_io_gpio_inst_GPIO61
		.hps_io_gpio_inst_GPIO65  (sys_hps_hps_io_hps_io_gpio_inst_GPIO65),                  //                  .hps_io_gpio_inst_GPIO65
		.h2f_rst_n                (sys_hps_h2f_reset_reset_n),                               //         h2f_reset.reset_n
		.f2h_sdram0_clk           (sys_hps_h2f_user1_clock_clk),                             //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_1_sys_hps_f2h_sdram0_data_address),       //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_1_sys_hps_f2h_sdram0_data_burstcount),    //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_1_sys_hps_f2h_sdram0_data_waitrequest),   //                  .waitrequest
		.f2h_sdram0_READDATA      (mm_interconnect_1_sys_hps_f2h_sdram0_data_readdata),      //                  .readdata
		.f2h_sdram0_READDATAVALID (mm_interconnect_1_sys_hps_f2h_sdram0_data_readdatavalid), //                  .readdatavalid
		.f2h_sdram0_READ          (mm_interconnect_1_sys_hps_f2h_sdram0_data_read),          //                  .read
		.f2h_sdram0_WRITEDATA     (mm_interconnect_1_sys_hps_f2h_sdram0_data_writedata),     //                  .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_1_sys_hps_f2h_sdram0_data_byteenable),    //                  .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_1_sys_hps_f2h_sdram0_data_write),         //                  .write
		.f2h_sdram1_clk           (sys_hps_h2f_user1_clock_clk),                             //  f2h_sdram1_clock.clk
		.f2h_sdram1_ARADDR        (),                                                        //   f2h_sdram1_data.araddr
		.f2h_sdram1_ARLEN         (),                                                        //                  .arlen
		.f2h_sdram1_ARID          (),                                                        //                  .arid
		.f2h_sdram1_ARSIZE        (),                                                        //                  .arsize
		.f2h_sdram1_ARBURST       (),                                                        //                  .arburst
		.f2h_sdram1_ARLOCK        (),                                                        //                  .arlock
		.f2h_sdram1_ARPROT        (),                                                        //                  .arprot
		.f2h_sdram1_ARVALID       (),                                                        //                  .arvalid
		.f2h_sdram1_ARCACHE       (),                                                        //                  .arcache
		.f2h_sdram1_AWADDR        (),                                                        //                  .awaddr
		.f2h_sdram1_AWLEN         (),                                                        //                  .awlen
		.f2h_sdram1_AWID          (),                                                        //                  .awid
		.f2h_sdram1_AWSIZE        (),                                                        //                  .awsize
		.f2h_sdram1_AWBURST       (),                                                        //                  .awburst
		.f2h_sdram1_AWLOCK        (),                                                        //                  .awlock
		.f2h_sdram1_AWPROT        (),                                                        //                  .awprot
		.f2h_sdram1_AWVALID       (),                                                        //                  .awvalid
		.f2h_sdram1_AWCACHE       (),                                                        //                  .awcache
		.f2h_sdram1_BRESP         (),                                                        //                  .bresp
		.f2h_sdram1_BID           (),                                                        //                  .bid
		.f2h_sdram1_BVALID        (),                                                        //                  .bvalid
		.f2h_sdram1_BREADY        (),                                                        //                  .bready
		.f2h_sdram1_ARREADY       (),                                                        //                  .arready
		.f2h_sdram1_AWREADY       (),                                                        //                  .awready
		.f2h_sdram1_RREADY        (),                                                        //                  .rready
		.f2h_sdram1_RDATA         (),                                                        //                  .rdata
		.f2h_sdram1_RRESP         (),                                                        //                  .rresp
		.f2h_sdram1_RLAST         (),                                                        //                  .rlast
		.f2h_sdram1_RID           (),                                                        //                  .rid
		.f2h_sdram1_RVALID        (),                                                        //                  .rvalid
		.f2h_sdram1_WLAST         (),                                                        //                  .wlast
		.f2h_sdram1_WVALID        (),                                                        //                  .wvalid
		.f2h_sdram1_WDATA         (),                                                        //                  .wdata
		.f2h_sdram1_WSTRB         (),                                                        //                  .wstrb
		.f2h_sdram1_WREADY        (),                                                        //                  .wready
		.f2h_sdram1_WID           (),                                                        //                  .wid
		.f2h_sdram2_clk           (sys_hps_h2f_user1_clock_clk),                             //  f2h_sdram2_clock.clk
		.f2h_sdram2_ARADDR        (),                                                        //   f2h_sdram2_data.araddr
		.f2h_sdram2_ARLEN         (),                                                        //                  .arlen
		.f2h_sdram2_ARID          (),                                                        //                  .arid
		.f2h_sdram2_ARSIZE        (),                                                        //                  .arsize
		.f2h_sdram2_ARBURST       (),                                                        //                  .arburst
		.f2h_sdram2_ARLOCK        (),                                                        //                  .arlock
		.f2h_sdram2_ARPROT        (),                                                        //                  .arprot
		.f2h_sdram2_ARVALID       (),                                                        //                  .arvalid
		.f2h_sdram2_ARCACHE       (),                                                        //                  .arcache
		.f2h_sdram2_AWADDR        (),                                                        //                  .awaddr
		.f2h_sdram2_AWLEN         (),                                                        //                  .awlen
		.f2h_sdram2_AWID          (),                                                        //                  .awid
		.f2h_sdram2_AWSIZE        (),                                                        //                  .awsize
		.f2h_sdram2_AWBURST       (),                                                        //                  .awburst
		.f2h_sdram2_AWLOCK        (),                                                        //                  .awlock
		.f2h_sdram2_AWPROT        (),                                                        //                  .awprot
		.f2h_sdram2_AWVALID       (),                                                        //                  .awvalid
		.f2h_sdram2_AWCACHE       (),                                                        //                  .awcache
		.f2h_sdram2_BRESP         (),                                                        //                  .bresp
		.f2h_sdram2_BID           (),                                                        //                  .bid
		.f2h_sdram2_BVALID        (),                                                        //                  .bvalid
		.f2h_sdram2_BREADY        (),                                                        //                  .bready
		.f2h_sdram2_ARREADY       (),                                                        //                  .arready
		.f2h_sdram2_AWREADY       (),                                                        //                  .awready
		.f2h_sdram2_RREADY        (),                                                        //                  .rready
		.f2h_sdram2_RDATA         (),                                                        //                  .rdata
		.f2h_sdram2_RRESP         (),                                                        //                  .rresp
		.f2h_sdram2_RLAST         (),                                                        //                  .rlast
		.f2h_sdram2_RID           (),                                                        //                  .rid
		.f2h_sdram2_RVALID        (),                                                        //                  .rvalid
		.f2h_sdram2_WLAST         (),                                                        //                  .wlast
		.f2h_sdram2_WVALID        (),                                                        //                  .wvalid
		.f2h_sdram2_WDATA         (),                                                        //                  .wdata
		.f2h_sdram2_WSTRB         (),                                                        //                  .wstrb
		.f2h_sdram2_WREADY        (),                                                        //                  .wready
		.f2h_sdram2_WID           (),                                                        //                  .wid
		.h2f_axi_clk              (sys_hps_h2f_user1_clock_clk),                             //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                                        //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                                        //                  .awaddr
		.h2f_AWLEN                (),                                                        //                  .awlen
		.h2f_AWSIZE               (),                                                        //                  .awsize
		.h2f_AWBURST              (),                                                        //                  .awburst
		.h2f_AWLOCK               (),                                                        //                  .awlock
		.h2f_AWCACHE              (),                                                        //                  .awcache
		.h2f_AWPROT               (),                                                        //                  .awprot
		.h2f_AWVALID              (),                                                        //                  .awvalid
		.h2f_AWREADY              (),                                                        //                  .awready
		.h2f_WID                  (),                                                        //                  .wid
		.h2f_WDATA                (),                                                        //                  .wdata
		.h2f_WSTRB                (),                                                        //                  .wstrb
		.h2f_WLAST                (),                                                        //                  .wlast
		.h2f_WVALID               (),                                                        //                  .wvalid
		.h2f_WREADY               (),                                                        //                  .wready
		.h2f_BID                  (),                                                        //                  .bid
		.h2f_BRESP                (),                                                        //                  .bresp
		.h2f_BVALID               (),                                                        //                  .bvalid
		.h2f_BREADY               (),                                                        //                  .bready
		.h2f_ARID                 (),                                                        //                  .arid
		.h2f_ARADDR               (),                                                        //                  .araddr
		.h2f_ARLEN                (),                                                        //                  .arlen
		.h2f_ARSIZE               (),                                                        //                  .arsize
		.h2f_ARBURST              (),                                                        //                  .arburst
		.h2f_ARLOCK               (),                                                        //                  .arlock
		.h2f_ARCACHE              (),                                                        //                  .arcache
		.h2f_ARPROT               (),                                                        //                  .arprot
		.h2f_ARVALID              (),                                                        //                  .arvalid
		.h2f_ARREADY              (),                                                        //                  .arready
		.h2f_RID                  (),                                                        //                  .rid
		.h2f_RDATA                (),                                                        //                  .rdata
		.h2f_RRESP                (),                                                        //                  .rresp
		.h2f_RLAST                (),                                                        //                  .rlast
		.h2f_RVALID               (),                                                        //                  .rvalid
		.h2f_RREADY               (),                                                        //                  .rready
		.f2h_axi_clk              (sys_hps_h2f_user1_clock_clk),                             //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                                        //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                                        //                  .awaddr
		.f2h_AWLEN                (),                                                        //                  .awlen
		.f2h_AWSIZE               (),                                                        //                  .awsize
		.f2h_AWBURST              (),                                                        //                  .awburst
		.f2h_AWLOCK               (),                                                        //                  .awlock
		.f2h_AWCACHE              (),                                                        //                  .awcache
		.f2h_AWPROT               (),                                                        //                  .awprot
		.f2h_AWVALID              (),                                                        //                  .awvalid
		.f2h_AWREADY              (),                                                        //                  .awready
		.f2h_AWUSER               (),                                                        //                  .awuser
		.f2h_WID                  (),                                                        //                  .wid
		.f2h_WDATA                (),                                                        //                  .wdata
		.f2h_WSTRB                (),                                                        //                  .wstrb
		.f2h_WLAST                (),                                                        //                  .wlast
		.f2h_WVALID               (),                                                        //                  .wvalid
		.f2h_WREADY               (),                                                        //                  .wready
		.f2h_BID                  (),                                                        //                  .bid
		.f2h_BRESP                (),                                                        //                  .bresp
		.f2h_BVALID               (),                                                        //                  .bvalid
		.f2h_BREADY               (),                                                        //                  .bready
		.f2h_ARID                 (),                                                        //                  .arid
		.f2h_ARADDR               (),                                                        //                  .araddr
		.f2h_ARLEN                (),                                                        //                  .arlen
		.f2h_ARSIZE               (),                                                        //                  .arsize
		.f2h_ARBURST              (),                                                        //                  .arburst
		.f2h_ARLOCK               (),                                                        //                  .arlock
		.f2h_ARCACHE              (),                                                        //                  .arcache
		.f2h_ARPROT               (),                                                        //                  .arprot
		.f2h_ARVALID              (),                                                        //                  .arvalid
		.f2h_ARREADY              (),                                                        //                  .arready
		.f2h_ARUSER               (),                                                        //                  .aruser
		.f2h_RID                  (),                                                        //                  .rid
		.f2h_RDATA                (),                                                        //                  .rdata
		.f2h_RRESP                (),                                                        //                  .rresp
		.f2h_RLAST                (),                                                        //                  .rlast
		.f2h_RVALID               (),                                                        //                  .rvalid
		.f2h_RREADY               (),                                                        //                  .rready
		.h2f_lw_axi_clk           (sys_hps_h2f_user1_clock_clk),                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (sys_hps_h2f_lw_axi_master_awid),                          // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (sys_hps_h2f_lw_axi_master_awaddr),                        //                  .awaddr
		.h2f_lw_AWLEN             (sys_hps_h2f_lw_axi_master_awlen),                         //                  .awlen
		.h2f_lw_AWSIZE            (sys_hps_h2f_lw_axi_master_awsize),                        //                  .awsize
		.h2f_lw_AWBURST           (sys_hps_h2f_lw_axi_master_awburst),                       //                  .awburst
		.h2f_lw_AWLOCK            (sys_hps_h2f_lw_axi_master_awlock),                        //                  .awlock
		.h2f_lw_AWCACHE           (sys_hps_h2f_lw_axi_master_awcache),                       //                  .awcache
		.h2f_lw_AWPROT            (sys_hps_h2f_lw_axi_master_awprot),                        //                  .awprot
		.h2f_lw_AWVALID           (sys_hps_h2f_lw_axi_master_awvalid),                       //                  .awvalid
		.h2f_lw_AWREADY           (sys_hps_h2f_lw_axi_master_awready),                       //                  .awready
		.h2f_lw_WID               (sys_hps_h2f_lw_axi_master_wid),                           //                  .wid
		.h2f_lw_WDATA             (sys_hps_h2f_lw_axi_master_wdata),                         //                  .wdata
		.h2f_lw_WSTRB             (sys_hps_h2f_lw_axi_master_wstrb),                         //                  .wstrb
		.h2f_lw_WLAST             (sys_hps_h2f_lw_axi_master_wlast),                         //                  .wlast
		.h2f_lw_WVALID            (sys_hps_h2f_lw_axi_master_wvalid),                        //                  .wvalid
		.h2f_lw_WREADY            (sys_hps_h2f_lw_axi_master_wready),                        //                  .wready
		.h2f_lw_BID               (sys_hps_h2f_lw_axi_master_bid),                           //                  .bid
		.h2f_lw_BRESP             (sys_hps_h2f_lw_axi_master_bresp),                         //                  .bresp
		.h2f_lw_BVALID            (sys_hps_h2f_lw_axi_master_bvalid),                        //                  .bvalid
		.h2f_lw_BREADY            (sys_hps_h2f_lw_axi_master_bready),                        //                  .bready
		.h2f_lw_ARID              (sys_hps_h2f_lw_axi_master_arid),                          //                  .arid
		.h2f_lw_ARADDR            (sys_hps_h2f_lw_axi_master_araddr),                        //                  .araddr
		.h2f_lw_ARLEN             (sys_hps_h2f_lw_axi_master_arlen),                         //                  .arlen
		.h2f_lw_ARSIZE            (sys_hps_h2f_lw_axi_master_arsize),                        //                  .arsize
		.h2f_lw_ARBURST           (sys_hps_h2f_lw_axi_master_arburst),                       //                  .arburst
		.h2f_lw_ARLOCK            (sys_hps_h2f_lw_axi_master_arlock),                        //                  .arlock
		.h2f_lw_ARCACHE           (sys_hps_h2f_lw_axi_master_arcache),                       //                  .arcache
		.h2f_lw_ARPROT            (sys_hps_h2f_lw_axi_master_arprot),                        //                  .arprot
		.h2f_lw_ARVALID           (sys_hps_h2f_lw_axi_master_arvalid),                       //                  .arvalid
		.h2f_lw_ARREADY           (sys_hps_h2f_lw_axi_master_arready),                       //                  .arready
		.h2f_lw_RID               (sys_hps_h2f_lw_axi_master_rid),                           //                  .rid
		.h2f_lw_RDATA             (sys_hps_h2f_lw_axi_master_rdata),                         //                  .rdata
		.h2f_lw_RRESP             (sys_hps_h2f_lw_axi_master_rresp),                         //                  .rresp
		.h2f_lw_RLAST             (sys_hps_h2f_lw_axi_master_rlast),                         //                  .rlast
		.h2f_lw_RVALID            (sys_hps_h2f_lw_axi_master_rvalid),                        //                  .rvalid
		.h2f_lw_RREADY            (sys_hps_h2f_lw_axi_master_rready),                        //                  .rready
		.f2h_irq_p0               (sys_hps_f2h_irq0_irq),                                    //          f2h_irq0.irq
		.f2h_irq_p1               (sys_hps_f2h_irq1_irq)                                     //          f2h_irq1.irq
	);

	system_bd_sys_id sys_id (
		.clock    (sys_hps_h2f_user1_clock_clk),                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	util_cpack2_impl #(
		.NUM_OF_CHANNELS     (4),
		.SAMPLES_PER_CHANNEL (1),
		.SAMPLE_DATA_WIDTH   (16)
	) util_adc_pack (
		.clk                     (sys_hps_h2f_user1_clock_clk),                                                                                                           //                        clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                        //                      reset.reset
		.packed_fifo_wr_en       (util_adc_pack_if_packed_fifo_wr_en_valid),                                                                                              //       if_packed_fifo_wr_en.valid
		.packed_fifo_wr_sync     (util_adc_pack_if_packed_fifo_wr_sync_sync),                                                                                             //     if_packed_fifo_wr_sync.sync
		.packed_fifo_wr_data     (util_adc_pack_if_packed_fifo_wr_data_data),                                                                                             //     if_packed_fifo_wr_data.data
		.packed_fifo_wr_overflow (axi_adc_dma_if_fifo_wr_overflow_ovf),                                                                                                   // if_packed_fifo_wr_overflow.ovf
		.fifo_wr_overflow        (util_adc_pack_if_fifo_wr_overflow_ovf),                                                                                                 //        if_fifo_wr_overflow.ovf
		.enable                  ({util_adc_wfifo_dout_3_enable,util_adc_wfifo_dout_2_enable,util_adc_wfifo_dout_1_enable,util_adc_wfifo_dout_0_enable}),                 //                   adc_ch_0.enable
		.fifo_wr_en              ({util_adc_wfifo_dout_3_valid,util_adc_wfifo_dout_2_valid,util_adc_wfifo_dout_1_valid,util_adc_wfifo_dout_0_valid}),                     //                           .valid
		.fifo_wr_data            ({util_adc_wfifo_dout_3_data[15:0],util_adc_wfifo_dout_2_data[15:0],util_adc_wfifo_dout_1_data[15:0],util_adc_wfifo_dout_0_data[15:0]})  //                           .data
	);

	util_wfifo #(
		.NUM_OF_CHANNELS   (4),
		.DIN_DATA_WIDTH    (16),
		.DOUT_DATA_WIDTH   (16),
		.DIN_ADDRESS_WIDTH (5)
	) util_adc_wfifo (
		.din_clk       (axi_adrv9001_if_adc_1_clk_clk),         //   if_din_clk.clk
		.din_rst       (axi_adrv9001_if_adc_1_rst_reset),       //   if_din_rst.reset
		.dout_clk      (sys_hps_h2f_user1_clock_clk),           //  if_dout_clk.clk
		.dout_rstn     (~rst_controller_reset_out_reset),       // if_dout_rstn.reset_n
		.din_enable_0  (axi_adrv9001_adc_1_ch_0_enable),        //        din_0.enable
		.din_valid_0   (axi_adrv9001_adc_1_ch_0_valid),         //             .valid
		.din_data_0    (axi_adrv9001_adc_1_ch_0_data),          //             .data
		.dout_enable_0 (util_adc_wfifo_dout_0_enable),          //       dout_0.enable
		.dout_valid_0  (util_adc_wfifo_dout_0_valid),           //             .valid
		.dout_data_0   (util_adc_wfifo_dout_0_data),            //             .data
		.din_ovf       (util_adc_wfifo_if_din_ovf_ovf),         //   if_din_ovf.ovf
		.dout_ovf      (util_adc_pack_if_fifo_wr_overflow_ovf), //  if_dout_ovf.ovf
		.din_enable_1  (axi_adrv9001_adc_1_ch_1_enable),        //        din_1.enable
		.din_valid_1   (axi_adrv9001_adc_1_ch_1_valid),         //             .valid
		.din_data_1    (axi_adrv9001_adc_1_ch_1_data),          //             .data
		.dout_enable_1 (util_adc_wfifo_dout_1_enable),          //       dout_1.enable
		.dout_valid_1  (util_adc_wfifo_dout_1_valid),           //             .valid
		.dout_data_1   (util_adc_wfifo_dout_1_data),            //             .data
		.din_enable_2  (axi_adrv9001_adc_1_ch_2_enable),        //        din_2.enable
		.din_valid_2   (axi_adrv9001_adc_1_ch_2_valid),         //             .valid
		.din_data_2    (axi_adrv9001_adc_1_ch_2_data),          //             .data
		.dout_enable_2 (util_adc_wfifo_dout_2_enable),          //       dout_2.enable
		.dout_valid_2  (util_adc_wfifo_dout_2_valid),           //             .valid
		.dout_data_2   (util_adc_wfifo_dout_2_data),            //             .data
		.din_enable_3  (axi_adrv9001_adc_1_ch_3_enable),        //        din_3.enable
		.din_valid_3   (axi_adrv9001_adc_1_ch_3_valid),         //             .valid
		.din_data_3    (axi_adrv9001_adc_1_ch_3_data),          //             .data
		.dout_enable_3 (util_adc_wfifo_dout_3_enable),          //       dout_3.enable
		.dout_valid_3  (util_adc_wfifo_dout_3_valid),           //             .valid
		.dout_data_3   (util_adc_wfifo_dout_3_data)             //             .data
	);

	util_rfifo #(
		.NUM_OF_CHANNELS   (4),
		.DIN_DATA_WIDTH    (16),
		.DOUT_DATA_WIDTH   (16),
		.DIN_ADDRESS_WIDTH (5)
	) util_dac_rfifo (
		.din_clk          (sys_hps_h2f_user1_clock_clk),             //  if_din_clk.clk
		.din_rstn         (~rst_controller_reset_out_reset),         // if_din_rstn.reset_n
		.dout_clk         (axi_adrv9001_if_dac_1_clk_clk),           // if_dout_clk.clk
		.dout_rst         (axi_adrv9001_if_dac_1_rst_reset),         // if_dout_rst.reset
		.din_enable_0     (util_dac_rfifo_din_0_enable),             //       din_0.enable
		.din_valid_0      (util_dac_rfifo_din_0_valid),              //            .valid
		.din_valid_in_0   (util_dac_upack_dac_ch_0_data_valid),      //            .data_valid
		.din_data_0       (util_dac_upack_dac_ch_0_data),            //            .data
		.dout_enable_0    (axi_adrv9001_dac_1_ch_0_enable),          //      dout_0.enable
		.dout_valid_0     (axi_adrv9001_dac_1_ch_0_valid),           //            .valid
		.dout_valid_out_0 (),                                        //            .data_valid
		.dout_data_0      (util_dac_rfifo_dout_0_data),              //            .data
		.din_unf          (util_dac_upack_if_fifo_rd_underflow_unf), //  if_din_unf.unf
		.dout_unf         (util_dac_rfifo_if_dout_unf_unf),          // if_dout_unf.unf
		.din_enable_1     (util_dac_rfifo_din_1_enable),             //       din_1.enable
		.din_valid_1      (util_dac_rfifo_din_1_valid),              //            .valid
		.din_valid_in_1   (util_dac_upack_dac_ch_1_data_valid),      //            .data_valid
		.din_data_1       (util_dac_upack_dac_ch_1_data),            //            .data
		.dout_enable_1    (axi_adrv9001_dac_1_ch_1_enable),          //      dout_1.enable
		.dout_valid_1     (axi_adrv9001_dac_1_ch_1_valid),           //            .valid
		.dout_valid_out_1 (),                                        //            .data_valid
		.dout_data_1      (util_dac_rfifo_dout_1_data),              //            .data
		.din_enable_2     (util_dac_rfifo_din_2_enable),             //       din_2.enable
		.din_valid_2      (util_dac_rfifo_din_2_valid),              //            .valid
		.din_valid_in_2   (util_dac_upack_dac_ch_2_data_valid),      //            .data_valid
		.din_data_2       (util_dac_upack_dac_ch_2_data),            //            .data
		.dout_enable_2    (axi_adrv9001_dac_1_ch_2_enable),          //      dout_2.enable
		.dout_valid_2     (axi_adrv9001_dac_1_ch_2_valid),           //            .valid
		.dout_valid_out_2 (),                                        //            .data_valid
		.dout_data_2      (util_dac_rfifo_dout_2_data),              //            .data
		.din_enable_3     (util_dac_rfifo_din_3_enable),             //       din_3.enable
		.din_valid_3      (util_dac_rfifo_din_3_valid),              //            .valid
		.din_valid_in_3   (util_dac_upack_dac_ch_3_data_valid),      //            .data_valid
		.din_data_3       (util_dac_upack_dac_ch_3_data),            //            .data
		.dout_enable_3    (axi_adrv9001_dac_1_ch_3_enable),          //      dout_3.enable
		.dout_valid_3     (axi_adrv9001_dac_1_ch_3_valid),           //            .valid
		.dout_valid_out_3 (),                                        //            .data_valid
		.dout_data_3      (util_dac_rfifo_dout_3_data)               //            .data
	);

	util_upack2_impl #(
		.NUM_OF_CHANNELS     (4),
		.SAMPLES_PER_CHANNEL (1),
		.SAMPLE_DATA_WIDTH   (16)
	) util_dac_upack (
		.clk               (sys_hps_h2f_user1_clock_clk),                                                                                                                  //                  clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                                                               //                reset.reset
		.s_axis_valid      (axi_dac_dma_m_axis_tvalid),                                                                                                                    //               s_axis.tvalid
		.s_axis_ready      (axi_dac_dma_m_axis_tready),                                                                                                                    //                     .tready
		.s_axis_data       (axi_dac_dma_m_axis_tdata),                                                                                                                     //                     .tdata
		.fifo_rd_underflow (util_dac_upack_if_fifo_rd_underflow_unf),                                                                                                      // if_fifo_rd_underflow.unf
		.enable            ({util_dac_rfifo_din_3_enable,util_dac_rfifo_din_2_enable,util_dac_rfifo_din_1_enable,util_dac_rfifo_din_0_enable}),                            //             dac_ch_0.enable
		.fifo_rd_en        ({util_dac_rfifo_din_3_valid,util_dac_rfifo_din_2_valid,util_dac_rfifo_din_1_valid,util_dac_rfifo_din_0_valid}),                                //                     .valid
		.fifo_rd_valid     (util_dac_upack_fifo_rd_valid[0]),                                                                                                              //                     .data_valid
		.fifo_rd_data      ({util_dac_upack_fifo_rd_data[63:48],util_dac_upack_fifo_rd_data[47:32],util_dac_upack_fifo_rd_data[31:16],util_dac_upack_fifo_rd_data[15:0]})  //                     .data
	);

	system_bd_mm_interconnect_0 mm_interconnect_0 (
		.axi_adc_dma_s_axi_awaddr                                              (mm_interconnect_0_axi_adc_dma_s_axi_awaddr),          //                                               axi_adc_dma_s_axi.awaddr
		.axi_adc_dma_s_axi_awprot                                              (mm_interconnect_0_axi_adc_dma_s_axi_awprot),          //                                                                .awprot
		.axi_adc_dma_s_axi_awvalid                                             (mm_interconnect_0_axi_adc_dma_s_axi_awvalid),         //                                                                .awvalid
		.axi_adc_dma_s_axi_awready                                             (mm_interconnect_0_axi_adc_dma_s_axi_awready),         //                                                                .awready
		.axi_adc_dma_s_axi_wdata                                               (mm_interconnect_0_axi_adc_dma_s_axi_wdata),           //                                                                .wdata
		.axi_adc_dma_s_axi_wstrb                                               (mm_interconnect_0_axi_adc_dma_s_axi_wstrb),           //                                                                .wstrb
		.axi_adc_dma_s_axi_wvalid                                              (mm_interconnect_0_axi_adc_dma_s_axi_wvalid),          //                                                                .wvalid
		.axi_adc_dma_s_axi_wready                                              (mm_interconnect_0_axi_adc_dma_s_axi_wready),          //                                                                .wready
		.axi_adc_dma_s_axi_bresp                                               (mm_interconnect_0_axi_adc_dma_s_axi_bresp),           //                                                                .bresp
		.axi_adc_dma_s_axi_bvalid                                              (mm_interconnect_0_axi_adc_dma_s_axi_bvalid),          //                                                                .bvalid
		.axi_adc_dma_s_axi_bready                                              (mm_interconnect_0_axi_adc_dma_s_axi_bready),          //                                                                .bready
		.axi_adc_dma_s_axi_araddr                                              (mm_interconnect_0_axi_adc_dma_s_axi_araddr),          //                                                                .araddr
		.axi_adc_dma_s_axi_arprot                                              (mm_interconnect_0_axi_adc_dma_s_axi_arprot),          //                                                                .arprot
		.axi_adc_dma_s_axi_arvalid                                             (mm_interconnect_0_axi_adc_dma_s_axi_arvalid),         //                                                                .arvalid
		.axi_adc_dma_s_axi_arready                                             (mm_interconnect_0_axi_adc_dma_s_axi_arready),         //                                                                .arready
		.axi_adc_dma_s_axi_rdata                                               (mm_interconnect_0_axi_adc_dma_s_axi_rdata),           //                                                                .rdata
		.axi_adc_dma_s_axi_rresp                                               (mm_interconnect_0_axi_adc_dma_s_axi_rresp),           //                                                                .rresp
		.axi_adc_dma_s_axi_rvalid                                              (mm_interconnect_0_axi_adc_dma_s_axi_rvalid),          //                                                                .rvalid
		.axi_adc_dma_s_axi_rready                                              (mm_interconnect_0_axi_adc_dma_s_axi_rready),          //                                                                .rready
		.axi_adrv9001_s_axi_awaddr                                             (mm_interconnect_0_axi_adrv9001_s_axi_awaddr),         //                                              axi_adrv9001_s_axi.awaddr
		.axi_adrv9001_s_axi_awprot                                             (mm_interconnect_0_axi_adrv9001_s_axi_awprot),         //                                                                .awprot
		.axi_adrv9001_s_axi_awvalid                                            (mm_interconnect_0_axi_adrv9001_s_axi_awvalid),        //                                                                .awvalid
		.axi_adrv9001_s_axi_awready                                            (mm_interconnect_0_axi_adrv9001_s_axi_awready),        //                                                                .awready
		.axi_adrv9001_s_axi_wdata                                              (mm_interconnect_0_axi_adrv9001_s_axi_wdata),          //                                                                .wdata
		.axi_adrv9001_s_axi_wstrb                                              (mm_interconnect_0_axi_adrv9001_s_axi_wstrb),          //                                                                .wstrb
		.axi_adrv9001_s_axi_wvalid                                             (mm_interconnect_0_axi_adrv9001_s_axi_wvalid),         //                                                                .wvalid
		.axi_adrv9001_s_axi_wready                                             (mm_interconnect_0_axi_adrv9001_s_axi_wready),         //                                                                .wready
		.axi_adrv9001_s_axi_bresp                                              (mm_interconnect_0_axi_adrv9001_s_axi_bresp),          //                                                                .bresp
		.axi_adrv9001_s_axi_bvalid                                             (mm_interconnect_0_axi_adrv9001_s_axi_bvalid),         //                                                                .bvalid
		.axi_adrv9001_s_axi_bready                                             (mm_interconnect_0_axi_adrv9001_s_axi_bready),         //                                                                .bready
		.axi_adrv9001_s_axi_araddr                                             (mm_interconnect_0_axi_adrv9001_s_axi_araddr),         //                                                                .araddr
		.axi_adrv9001_s_axi_arprot                                             (mm_interconnect_0_axi_adrv9001_s_axi_arprot),         //                                                                .arprot
		.axi_adrv9001_s_axi_arvalid                                            (mm_interconnect_0_axi_adrv9001_s_axi_arvalid),        //                                                                .arvalid
		.axi_adrv9001_s_axi_arready                                            (mm_interconnect_0_axi_adrv9001_s_axi_arready),        //                                                                .arready
		.axi_adrv9001_s_axi_rdata                                              (mm_interconnect_0_axi_adrv9001_s_axi_rdata),          //                                                                .rdata
		.axi_adrv9001_s_axi_rresp                                              (mm_interconnect_0_axi_adrv9001_s_axi_rresp),          //                                                                .rresp
		.axi_adrv9001_s_axi_rvalid                                             (mm_interconnect_0_axi_adrv9001_s_axi_rvalid),         //                                                                .rvalid
		.axi_adrv9001_s_axi_rready                                             (mm_interconnect_0_axi_adrv9001_s_axi_rready),         //                                                                .rready
		.axi_dac_dma_s_axi_awaddr                                              (mm_interconnect_0_axi_dac_dma_s_axi_awaddr),          //                                               axi_dac_dma_s_axi.awaddr
		.axi_dac_dma_s_axi_awprot                                              (mm_interconnect_0_axi_dac_dma_s_axi_awprot),          //                                                                .awprot
		.axi_dac_dma_s_axi_awvalid                                             (mm_interconnect_0_axi_dac_dma_s_axi_awvalid),         //                                                                .awvalid
		.axi_dac_dma_s_axi_awready                                             (mm_interconnect_0_axi_dac_dma_s_axi_awready),         //                                                                .awready
		.axi_dac_dma_s_axi_wdata                                               (mm_interconnect_0_axi_dac_dma_s_axi_wdata),           //                                                                .wdata
		.axi_dac_dma_s_axi_wstrb                                               (mm_interconnect_0_axi_dac_dma_s_axi_wstrb),           //                                                                .wstrb
		.axi_dac_dma_s_axi_wvalid                                              (mm_interconnect_0_axi_dac_dma_s_axi_wvalid),          //                                                                .wvalid
		.axi_dac_dma_s_axi_wready                                              (mm_interconnect_0_axi_dac_dma_s_axi_wready),          //                                                                .wready
		.axi_dac_dma_s_axi_bresp                                               (mm_interconnect_0_axi_dac_dma_s_axi_bresp),           //                                                                .bresp
		.axi_dac_dma_s_axi_bvalid                                              (mm_interconnect_0_axi_dac_dma_s_axi_bvalid),          //                                                                .bvalid
		.axi_dac_dma_s_axi_bready                                              (mm_interconnect_0_axi_dac_dma_s_axi_bready),          //                                                                .bready
		.axi_dac_dma_s_axi_araddr                                              (mm_interconnect_0_axi_dac_dma_s_axi_araddr),          //                                                                .araddr
		.axi_dac_dma_s_axi_arprot                                              (mm_interconnect_0_axi_dac_dma_s_axi_arprot),          //                                                                .arprot
		.axi_dac_dma_s_axi_arvalid                                             (mm_interconnect_0_axi_dac_dma_s_axi_arvalid),         //                                                                .arvalid
		.axi_dac_dma_s_axi_arready                                             (mm_interconnect_0_axi_dac_dma_s_axi_arready),         //                                                                .arready
		.axi_dac_dma_s_axi_rdata                                               (mm_interconnect_0_axi_dac_dma_s_axi_rdata),           //                                                                .rdata
		.axi_dac_dma_s_axi_rresp                                               (mm_interconnect_0_axi_dac_dma_s_axi_rresp),           //                                                                .rresp
		.axi_dac_dma_s_axi_rvalid                                              (mm_interconnect_0_axi_dac_dma_s_axi_rvalid),          //                                                                .rvalid
		.axi_dac_dma_s_axi_rready                                              (mm_interconnect_0_axi_dac_dma_s_axi_rready),          //                                                                .rready
		.axi_hdmi_tx_0_s_axi_awaddr                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awaddr),        //                                             axi_hdmi_tx_0_s_axi.awaddr
		.axi_hdmi_tx_0_s_axi_awprot                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awprot),        //                                                                .awprot
		.axi_hdmi_tx_0_s_axi_awvalid                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awvalid),       //                                                                .awvalid
		.axi_hdmi_tx_0_s_axi_awready                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_awready),       //                                                                .awready
		.axi_hdmi_tx_0_s_axi_wdata                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wdata),         //                                                                .wdata
		.axi_hdmi_tx_0_s_axi_wstrb                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wstrb),         //                                                                .wstrb
		.axi_hdmi_tx_0_s_axi_wvalid                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wvalid),        //                                                                .wvalid
		.axi_hdmi_tx_0_s_axi_wready                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_wready),        //                                                                .wready
		.axi_hdmi_tx_0_s_axi_bresp                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bresp),         //                                                                .bresp
		.axi_hdmi_tx_0_s_axi_bvalid                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bvalid),        //                                                                .bvalid
		.axi_hdmi_tx_0_s_axi_bready                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_bready),        //                                                                .bready
		.axi_hdmi_tx_0_s_axi_araddr                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_araddr),        //                                                                .araddr
		.axi_hdmi_tx_0_s_axi_arprot                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arprot),        //                                                                .arprot
		.axi_hdmi_tx_0_s_axi_arvalid                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arvalid),       //                                                                .arvalid
		.axi_hdmi_tx_0_s_axi_arready                                           (mm_interconnect_0_axi_hdmi_tx_0_s_axi_arready),       //                                                                .arready
		.axi_hdmi_tx_0_s_axi_rdata                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rdata),         //                                                                .rdata
		.axi_hdmi_tx_0_s_axi_rresp                                             (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rresp),         //                                                                .rresp
		.axi_hdmi_tx_0_s_axi_rvalid                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rvalid),        //                                                                .rvalid
		.axi_hdmi_tx_0_s_axi_rready                                            (mm_interconnect_0_axi_hdmi_tx_0_s_axi_rready),        //                                                                .rready
		.hdmi_dmac_0_s_axi_awaddr                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_awaddr),          //                                               hdmi_dmac_0_s_axi.awaddr
		.hdmi_dmac_0_s_axi_awprot                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_awprot),          //                                                                .awprot
		.hdmi_dmac_0_s_axi_awvalid                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_awvalid),         //                                                                .awvalid
		.hdmi_dmac_0_s_axi_awready                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_awready),         //                                                                .awready
		.hdmi_dmac_0_s_axi_wdata                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_wdata),           //                                                                .wdata
		.hdmi_dmac_0_s_axi_wstrb                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_wstrb),           //                                                                .wstrb
		.hdmi_dmac_0_s_axi_wvalid                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_wvalid),          //                                                                .wvalid
		.hdmi_dmac_0_s_axi_wready                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_wready),          //                                                                .wready
		.hdmi_dmac_0_s_axi_bresp                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_bresp),           //                                                                .bresp
		.hdmi_dmac_0_s_axi_bvalid                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_bvalid),          //                                                                .bvalid
		.hdmi_dmac_0_s_axi_bready                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_bready),          //                                                                .bready
		.hdmi_dmac_0_s_axi_araddr                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_araddr),          //                                                                .araddr
		.hdmi_dmac_0_s_axi_arprot                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_arprot),          //                                                                .arprot
		.hdmi_dmac_0_s_axi_arvalid                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_arvalid),         //                                                                .arvalid
		.hdmi_dmac_0_s_axi_arready                                             (mm_interconnect_0_hdmi_dmac_0_s_axi_arready),         //                                                                .arready
		.hdmi_dmac_0_s_axi_rdata                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_rdata),           //                                                                .rdata
		.hdmi_dmac_0_s_axi_rresp                                               (mm_interconnect_0_hdmi_dmac_0_s_axi_rresp),           //                                                                .rresp
		.hdmi_dmac_0_s_axi_rvalid                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_rvalid),          //                                                                .rvalid
		.hdmi_dmac_0_s_axi_rready                                              (mm_interconnect_0_hdmi_dmac_0_s_axi_rready),          //                                                                .rready
		.sys_hps_h2f_lw_axi_master_awid                                        (sys_hps_h2f_lw_axi_master_awid),                      //                                       sys_hps_h2f_lw_axi_master.awid
		.sys_hps_h2f_lw_axi_master_awaddr                                      (sys_hps_h2f_lw_axi_master_awaddr),                    //                                                                .awaddr
		.sys_hps_h2f_lw_axi_master_awlen                                       (sys_hps_h2f_lw_axi_master_awlen),                     //                                                                .awlen
		.sys_hps_h2f_lw_axi_master_awsize                                      (sys_hps_h2f_lw_axi_master_awsize),                    //                                                                .awsize
		.sys_hps_h2f_lw_axi_master_awburst                                     (sys_hps_h2f_lw_axi_master_awburst),                   //                                                                .awburst
		.sys_hps_h2f_lw_axi_master_awlock                                      (sys_hps_h2f_lw_axi_master_awlock),                    //                                                                .awlock
		.sys_hps_h2f_lw_axi_master_awcache                                     (sys_hps_h2f_lw_axi_master_awcache),                   //                                                                .awcache
		.sys_hps_h2f_lw_axi_master_awprot                                      (sys_hps_h2f_lw_axi_master_awprot),                    //                                                                .awprot
		.sys_hps_h2f_lw_axi_master_awvalid                                     (sys_hps_h2f_lw_axi_master_awvalid),                   //                                                                .awvalid
		.sys_hps_h2f_lw_axi_master_awready                                     (sys_hps_h2f_lw_axi_master_awready),                   //                                                                .awready
		.sys_hps_h2f_lw_axi_master_wid                                         (sys_hps_h2f_lw_axi_master_wid),                       //                                                                .wid
		.sys_hps_h2f_lw_axi_master_wdata                                       (sys_hps_h2f_lw_axi_master_wdata),                     //                                                                .wdata
		.sys_hps_h2f_lw_axi_master_wstrb                                       (sys_hps_h2f_lw_axi_master_wstrb),                     //                                                                .wstrb
		.sys_hps_h2f_lw_axi_master_wlast                                       (sys_hps_h2f_lw_axi_master_wlast),                     //                                                                .wlast
		.sys_hps_h2f_lw_axi_master_wvalid                                      (sys_hps_h2f_lw_axi_master_wvalid),                    //                                                                .wvalid
		.sys_hps_h2f_lw_axi_master_wready                                      (sys_hps_h2f_lw_axi_master_wready),                    //                                                                .wready
		.sys_hps_h2f_lw_axi_master_bid                                         (sys_hps_h2f_lw_axi_master_bid),                       //                                                                .bid
		.sys_hps_h2f_lw_axi_master_bresp                                       (sys_hps_h2f_lw_axi_master_bresp),                     //                                                                .bresp
		.sys_hps_h2f_lw_axi_master_bvalid                                      (sys_hps_h2f_lw_axi_master_bvalid),                    //                                                                .bvalid
		.sys_hps_h2f_lw_axi_master_bready                                      (sys_hps_h2f_lw_axi_master_bready),                    //                                                                .bready
		.sys_hps_h2f_lw_axi_master_arid                                        (sys_hps_h2f_lw_axi_master_arid),                      //                                                                .arid
		.sys_hps_h2f_lw_axi_master_araddr                                      (sys_hps_h2f_lw_axi_master_araddr),                    //                                                                .araddr
		.sys_hps_h2f_lw_axi_master_arlen                                       (sys_hps_h2f_lw_axi_master_arlen),                     //                                                                .arlen
		.sys_hps_h2f_lw_axi_master_arsize                                      (sys_hps_h2f_lw_axi_master_arsize),                    //                                                                .arsize
		.sys_hps_h2f_lw_axi_master_arburst                                     (sys_hps_h2f_lw_axi_master_arburst),                   //                                                                .arburst
		.sys_hps_h2f_lw_axi_master_arlock                                      (sys_hps_h2f_lw_axi_master_arlock),                    //                                                                .arlock
		.sys_hps_h2f_lw_axi_master_arcache                                     (sys_hps_h2f_lw_axi_master_arcache),                   //                                                                .arcache
		.sys_hps_h2f_lw_axi_master_arprot                                      (sys_hps_h2f_lw_axi_master_arprot),                    //                                                                .arprot
		.sys_hps_h2f_lw_axi_master_arvalid                                     (sys_hps_h2f_lw_axi_master_arvalid),                   //                                                                .arvalid
		.sys_hps_h2f_lw_axi_master_arready                                     (sys_hps_h2f_lw_axi_master_arready),                   //                                                                .arready
		.sys_hps_h2f_lw_axi_master_rid                                         (sys_hps_h2f_lw_axi_master_rid),                       //                                                                .rid
		.sys_hps_h2f_lw_axi_master_rdata                                       (sys_hps_h2f_lw_axi_master_rdata),                     //                                                                .rdata
		.sys_hps_h2f_lw_axi_master_rresp                                       (sys_hps_h2f_lw_axi_master_rresp),                     //                                                                .rresp
		.sys_hps_h2f_lw_axi_master_rlast                                       (sys_hps_h2f_lw_axi_master_rlast),                     //                                                                .rlast
		.sys_hps_h2f_lw_axi_master_rvalid                                      (sys_hps_h2f_lw_axi_master_rvalid),                    //                                                                .rvalid
		.sys_hps_h2f_lw_axi_master_rready                                      (sys_hps_h2f_lw_axi_master_rready),                    //                                                                .rready
		.sys_hps_h2f_user1_clock_clk                                           (sys_hps_h2f_user1_clock_clk),                         //                                         sys_hps_h2f_user1_clock.clk
		.sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // sys_hps_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.sys_id_reset_reset_bridge_in_reset_reset                              (rst_controller_reset_out_reset),                      //                              sys_id_reset_reset_bridge_in_reset.reset
		.avl_adrv9001_gpio_s1_address                                          (mm_interconnect_0_avl_adrv9001_gpio_s1_address),      //                                            avl_adrv9001_gpio_s1.address
		.avl_adrv9001_gpio_s1_write                                            (mm_interconnect_0_avl_adrv9001_gpio_s1_write),        //                                                                .write
		.avl_adrv9001_gpio_s1_readdata                                         (mm_interconnect_0_avl_adrv9001_gpio_s1_readdata),     //                                                                .readdata
		.avl_adrv9001_gpio_s1_writedata                                        (mm_interconnect_0_avl_adrv9001_gpio_s1_writedata),    //                                                                .writedata
		.avl_adrv9001_gpio_s1_chipselect                                       (mm_interconnect_0_avl_adrv9001_gpio_s1_chipselect),   //                                                                .chipselect
		.spi_0_spi_control_port_address                                        (mm_interconnect_0_spi_0_spi_control_port_address),    //                                          spi_0_spi_control_port.address
		.spi_0_spi_control_port_write                                          (mm_interconnect_0_spi_0_spi_control_port_write),      //                                                                .write
		.spi_0_spi_control_port_read                                           (mm_interconnect_0_spi_0_spi_control_port_read),       //                                                                .read
		.spi_0_spi_control_port_readdata                                       (mm_interconnect_0_spi_0_spi_control_port_readdata),   //                                                                .readdata
		.spi_0_spi_control_port_writedata                                      (mm_interconnect_0_spi_0_spi_control_port_writedata),  //                                                                .writedata
		.spi_0_spi_control_port_chipselect                                     (mm_interconnect_0_spi_0_spi_control_port_chipselect), //                                                                .chipselect
		.sys_gpio_bd_s1_address                                                (mm_interconnect_0_sys_gpio_bd_s1_address),            //                                                  sys_gpio_bd_s1.address
		.sys_gpio_bd_s1_write                                                  (mm_interconnect_0_sys_gpio_bd_s1_write),              //                                                                .write
		.sys_gpio_bd_s1_readdata                                               (mm_interconnect_0_sys_gpio_bd_s1_readdata),           //                                                                .readdata
		.sys_gpio_bd_s1_writedata                                              (mm_interconnect_0_sys_gpio_bd_s1_writedata),          //                                                                .writedata
		.sys_gpio_bd_s1_chipselect                                             (mm_interconnect_0_sys_gpio_bd_s1_chipselect),         //                                                                .chipselect
		.sys_gpio_in_s1_address                                                (mm_interconnect_0_sys_gpio_in_s1_address),            //                                                  sys_gpio_in_s1.address
		.sys_gpio_in_s1_write                                                  (mm_interconnect_0_sys_gpio_in_s1_write),              //                                                                .write
		.sys_gpio_in_s1_readdata                                               (mm_interconnect_0_sys_gpio_in_s1_readdata),           //                                                                .readdata
		.sys_gpio_in_s1_writedata                                              (mm_interconnect_0_sys_gpio_in_s1_writedata),          //                                                                .writedata
		.sys_gpio_in_s1_chipselect                                             (mm_interconnect_0_sys_gpio_in_s1_chipselect),         //                                                                .chipselect
		.sys_gpio_out_s1_address                                               (mm_interconnect_0_sys_gpio_out_s1_address),           //                                                 sys_gpio_out_s1.address
		.sys_gpio_out_s1_write                                                 (mm_interconnect_0_sys_gpio_out_s1_write),             //                                                                .write
		.sys_gpio_out_s1_readdata                                              (mm_interconnect_0_sys_gpio_out_s1_readdata),          //                                                                .readdata
		.sys_gpio_out_s1_writedata                                             (mm_interconnect_0_sys_gpio_out_s1_writedata),         //                                                                .writedata
		.sys_gpio_out_s1_chipselect                                            (mm_interconnect_0_sys_gpio_out_s1_chipselect),        //                                                                .chipselect
		.sys_id_control_slave_address                                          (mm_interconnect_0_sys_id_control_slave_address),      //                                            sys_id_control_slave.address
		.sys_id_control_slave_readdata                                         (mm_interconnect_0_sys_id_control_slave_readdata)      //                                                                .readdata
	);

	system_bd_mm_interconnect_1 mm_interconnect_1 (
		.axi_adc_dma_m_dest_axi_awid                                          (axi_adc_dma_m_dest_axi_awid),                             //                                         axi_adc_dma_m_dest_axi.awid
		.axi_adc_dma_m_dest_axi_awaddr                                        (axi_adc_dma_m_dest_axi_awaddr),                           //                                                               .awaddr
		.axi_adc_dma_m_dest_axi_awlen                                         (axi_adc_dma_m_dest_axi_awlen),                            //                                                               .awlen
		.axi_adc_dma_m_dest_axi_awsize                                        (axi_adc_dma_m_dest_axi_awsize),                           //                                                               .awsize
		.axi_adc_dma_m_dest_axi_awburst                                       (axi_adc_dma_m_dest_axi_awburst),                          //                                                               .awburst
		.axi_adc_dma_m_dest_axi_awlock                                        (axi_adc_dma_m_dest_axi_awlock),                           //                                                               .awlock
		.axi_adc_dma_m_dest_axi_awcache                                       (axi_adc_dma_m_dest_axi_awcache),                          //                                                               .awcache
		.axi_adc_dma_m_dest_axi_awprot                                        (axi_adc_dma_m_dest_axi_awprot),                           //                                                               .awprot
		.axi_adc_dma_m_dest_axi_awvalid                                       (axi_adc_dma_m_dest_axi_awvalid),                          //                                                               .awvalid
		.axi_adc_dma_m_dest_axi_awready                                       (axi_adc_dma_m_dest_axi_awready),                          //                                                               .awready
		.axi_adc_dma_m_dest_axi_wid                                           (axi_adc_dma_m_dest_axi_wid),                              //                                                               .wid
		.axi_adc_dma_m_dest_axi_wdata                                         (axi_adc_dma_m_dest_axi_wdata),                            //                                                               .wdata
		.axi_adc_dma_m_dest_axi_wstrb                                         (axi_adc_dma_m_dest_axi_wstrb),                            //                                                               .wstrb
		.axi_adc_dma_m_dest_axi_wlast                                         (axi_adc_dma_m_dest_axi_wlast),                            //                                                               .wlast
		.axi_adc_dma_m_dest_axi_wvalid                                        (axi_adc_dma_m_dest_axi_wvalid),                           //                                                               .wvalid
		.axi_adc_dma_m_dest_axi_wready                                        (axi_adc_dma_m_dest_axi_wready),                           //                                                               .wready
		.axi_adc_dma_m_dest_axi_bid                                           (axi_adc_dma_m_dest_axi_bid),                              //                                                               .bid
		.axi_adc_dma_m_dest_axi_bresp                                         (axi_adc_dma_m_dest_axi_bresp),                            //                                                               .bresp
		.axi_adc_dma_m_dest_axi_bvalid                                        (axi_adc_dma_m_dest_axi_bvalid),                           //                                                               .bvalid
		.axi_adc_dma_m_dest_axi_bready                                        (axi_adc_dma_m_dest_axi_bready),                           //                                                               .bready
		.axi_adc_dma_m_dest_axi_arid                                          (axi_adc_dma_m_dest_axi_arid),                             //                                                               .arid
		.axi_adc_dma_m_dest_axi_araddr                                        (axi_adc_dma_m_dest_axi_araddr),                           //                                                               .araddr
		.axi_adc_dma_m_dest_axi_arlen                                         (axi_adc_dma_m_dest_axi_arlen),                            //                                                               .arlen
		.axi_adc_dma_m_dest_axi_arsize                                        (axi_adc_dma_m_dest_axi_arsize),                           //                                                               .arsize
		.axi_adc_dma_m_dest_axi_arburst                                       (axi_adc_dma_m_dest_axi_arburst),                          //                                                               .arburst
		.axi_adc_dma_m_dest_axi_arlock                                        (axi_adc_dma_m_dest_axi_arlock),                           //                                                               .arlock
		.axi_adc_dma_m_dest_axi_arcache                                       (axi_adc_dma_m_dest_axi_arcache),                          //                                                               .arcache
		.axi_adc_dma_m_dest_axi_arprot                                        (axi_adc_dma_m_dest_axi_arprot),                           //                                                               .arprot
		.axi_adc_dma_m_dest_axi_arvalid                                       (axi_adc_dma_m_dest_axi_arvalid),                          //                                                               .arvalid
		.axi_adc_dma_m_dest_axi_arready                                       (axi_adc_dma_m_dest_axi_arready),                          //                                                               .arready
		.axi_adc_dma_m_dest_axi_rid                                           (axi_adc_dma_m_dest_axi_rid),                              //                                                               .rid
		.axi_adc_dma_m_dest_axi_rdata                                         (axi_adc_dma_m_dest_axi_rdata),                            //                                                               .rdata
		.axi_adc_dma_m_dest_axi_rresp                                         (axi_adc_dma_m_dest_axi_rresp),                            //                                                               .rresp
		.axi_adc_dma_m_dest_axi_rlast                                         (axi_adc_dma_m_dest_axi_rlast),                            //                                                               .rlast
		.axi_adc_dma_m_dest_axi_rvalid                                        (axi_adc_dma_m_dest_axi_rvalid),                           //                                                               .rvalid
		.axi_adc_dma_m_dest_axi_rready                                        (axi_adc_dma_m_dest_axi_rready),                           //                                                               .rready
		.axi_dac_dma_m_src_axi_awid                                           (axi_dac_dma_m_src_axi_awid),                              //                                          axi_dac_dma_m_src_axi.awid
		.axi_dac_dma_m_src_axi_awaddr                                         (axi_dac_dma_m_src_axi_awaddr),                            //                                                               .awaddr
		.axi_dac_dma_m_src_axi_awlen                                          (axi_dac_dma_m_src_axi_awlen),                             //                                                               .awlen
		.axi_dac_dma_m_src_axi_awsize                                         (axi_dac_dma_m_src_axi_awsize),                            //                                                               .awsize
		.axi_dac_dma_m_src_axi_awburst                                        (axi_dac_dma_m_src_axi_awburst),                           //                                                               .awburst
		.axi_dac_dma_m_src_axi_awlock                                         (axi_dac_dma_m_src_axi_awlock),                            //                                                               .awlock
		.axi_dac_dma_m_src_axi_awcache                                        (axi_dac_dma_m_src_axi_awcache),                           //                                                               .awcache
		.axi_dac_dma_m_src_axi_awprot                                         (axi_dac_dma_m_src_axi_awprot),                            //                                                               .awprot
		.axi_dac_dma_m_src_axi_awvalid                                        (axi_dac_dma_m_src_axi_awvalid),                           //                                                               .awvalid
		.axi_dac_dma_m_src_axi_awready                                        (axi_dac_dma_m_src_axi_awready),                           //                                                               .awready
		.axi_dac_dma_m_src_axi_wid                                            (axi_dac_dma_m_src_axi_wid),                               //                                                               .wid
		.axi_dac_dma_m_src_axi_wdata                                          (axi_dac_dma_m_src_axi_wdata),                             //                                                               .wdata
		.axi_dac_dma_m_src_axi_wstrb                                          (axi_dac_dma_m_src_axi_wstrb),                             //                                                               .wstrb
		.axi_dac_dma_m_src_axi_wlast                                          (axi_dac_dma_m_src_axi_wlast),                             //                                                               .wlast
		.axi_dac_dma_m_src_axi_wvalid                                         (axi_dac_dma_m_src_axi_wvalid),                            //                                                               .wvalid
		.axi_dac_dma_m_src_axi_wready                                         (axi_dac_dma_m_src_axi_wready),                            //                                                               .wready
		.axi_dac_dma_m_src_axi_bid                                            (axi_dac_dma_m_src_axi_bid),                               //                                                               .bid
		.axi_dac_dma_m_src_axi_bresp                                          (axi_dac_dma_m_src_axi_bresp),                             //                                                               .bresp
		.axi_dac_dma_m_src_axi_bvalid                                         (axi_dac_dma_m_src_axi_bvalid),                            //                                                               .bvalid
		.axi_dac_dma_m_src_axi_bready                                         (axi_dac_dma_m_src_axi_bready),                            //                                                               .bready
		.axi_dac_dma_m_src_axi_arid                                           (axi_dac_dma_m_src_axi_arid),                              //                                                               .arid
		.axi_dac_dma_m_src_axi_araddr                                         (axi_dac_dma_m_src_axi_araddr),                            //                                                               .araddr
		.axi_dac_dma_m_src_axi_arlen                                          (axi_dac_dma_m_src_axi_arlen),                             //                                                               .arlen
		.axi_dac_dma_m_src_axi_arsize                                         (axi_dac_dma_m_src_axi_arsize),                            //                                                               .arsize
		.axi_dac_dma_m_src_axi_arburst                                        (axi_dac_dma_m_src_axi_arburst),                           //                                                               .arburst
		.axi_dac_dma_m_src_axi_arlock                                         (axi_dac_dma_m_src_axi_arlock),                            //                                                               .arlock
		.axi_dac_dma_m_src_axi_arcache                                        (axi_dac_dma_m_src_axi_arcache),                           //                                                               .arcache
		.axi_dac_dma_m_src_axi_arprot                                         (axi_dac_dma_m_src_axi_arprot),                            //                                                               .arprot
		.axi_dac_dma_m_src_axi_arvalid                                        (axi_dac_dma_m_src_axi_arvalid),                           //                                                               .arvalid
		.axi_dac_dma_m_src_axi_arready                                        (axi_dac_dma_m_src_axi_arready),                           //                                                               .arready
		.axi_dac_dma_m_src_axi_rid                                            (axi_dac_dma_m_src_axi_rid),                               //                                                               .rid
		.axi_dac_dma_m_src_axi_rdata                                          (axi_dac_dma_m_src_axi_rdata),                             //                                                               .rdata
		.axi_dac_dma_m_src_axi_rresp                                          (axi_dac_dma_m_src_axi_rresp),                             //                                                               .rresp
		.axi_dac_dma_m_src_axi_rlast                                          (axi_dac_dma_m_src_axi_rlast),                             //                                                               .rlast
		.axi_dac_dma_m_src_axi_rvalid                                         (axi_dac_dma_m_src_axi_rvalid),                            //                                                               .rvalid
		.axi_dac_dma_m_src_axi_rready                                         (axi_dac_dma_m_src_axi_rready),                            //                                                               .rready
		.hdmi_dmac_0_m_src_axi_awid                                           (hdmi_dmac_0_m_src_axi_awid),                              //                                          hdmi_dmac_0_m_src_axi.awid
		.hdmi_dmac_0_m_src_axi_awaddr                                         (hdmi_dmac_0_m_src_axi_awaddr),                            //                                                               .awaddr
		.hdmi_dmac_0_m_src_axi_awlen                                          (hdmi_dmac_0_m_src_axi_awlen),                             //                                                               .awlen
		.hdmi_dmac_0_m_src_axi_awsize                                         (hdmi_dmac_0_m_src_axi_awsize),                            //                                                               .awsize
		.hdmi_dmac_0_m_src_axi_awburst                                        (hdmi_dmac_0_m_src_axi_awburst),                           //                                                               .awburst
		.hdmi_dmac_0_m_src_axi_awlock                                         (hdmi_dmac_0_m_src_axi_awlock),                            //                                                               .awlock
		.hdmi_dmac_0_m_src_axi_awcache                                        (hdmi_dmac_0_m_src_axi_awcache),                           //                                                               .awcache
		.hdmi_dmac_0_m_src_axi_awprot                                         (hdmi_dmac_0_m_src_axi_awprot),                            //                                                               .awprot
		.hdmi_dmac_0_m_src_axi_awvalid                                        (hdmi_dmac_0_m_src_axi_awvalid),                           //                                                               .awvalid
		.hdmi_dmac_0_m_src_axi_awready                                        (hdmi_dmac_0_m_src_axi_awready),                           //                                                               .awready
		.hdmi_dmac_0_m_src_axi_wid                                            (hdmi_dmac_0_m_src_axi_wid),                               //                                                               .wid
		.hdmi_dmac_0_m_src_axi_wdata                                          (hdmi_dmac_0_m_src_axi_wdata),                             //                                                               .wdata
		.hdmi_dmac_0_m_src_axi_wstrb                                          (hdmi_dmac_0_m_src_axi_wstrb),                             //                                                               .wstrb
		.hdmi_dmac_0_m_src_axi_wlast                                          (hdmi_dmac_0_m_src_axi_wlast),                             //                                                               .wlast
		.hdmi_dmac_0_m_src_axi_wvalid                                         (hdmi_dmac_0_m_src_axi_wvalid),                            //                                                               .wvalid
		.hdmi_dmac_0_m_src_axi_wready                                         (hdmi_dmac_0_m_src_axi_wready),                            //                                                               .wready
		.hdmi_dmac_0_m_src_axi_bid                                            (hdmi_dmac_0_m_src_axi_bid),                               //                                                               .bid
		.hdmi_dmac_0_m_src_axi_bresp                                          (hdmi_dmac_0_m_src_axi_bresp),                             //                                                               .bresp
		.hdmi_dmac_0_m_src_axi_bvalid                                         (hdmi_dmac_0_m_src_axi_bvalid),                            //                                                               .bvalid
		.hdmi_dmac_0_m_src_axi_bready                                         (hdmi_dmac_0_m_src_axi_bready),                            //                                                               .bready
		.hdmi_dmac_0_m_src_axi_arid                                           (hdmi_dmac_0_m_src_axi_arid),                              //                                                               .arid
		.hdmi_dmac_0_m_src_axi_araddr                                         (hdmi_dmac_0_m_src_axi_araddr),                            //                                                               .araddr
		.hdmi_dmac_0_m_src_axi_arlen                                          (hdmi_dmac_0_m_src_axi_arlen),                             //                                                               .arlen
		.hdmi_dmac_0_m_src_axi_arsize                                         (hdmi_dmac_0_m_src_axi_arsize),                            //                                                               .arsize
		.hdmi_dmac_0_m_src_axi_arburst                                        (hdmi_dmac_0_m_src_axi_arburst),                           //                                                               .arburst
		.hdmi_dmac_0_m_src_axi_arlock                                         (hdmi_dmac_0_m_src_axi_arlock),                            //                                                               .arlock
		.hdmi_dmac_0_m_src_axi_arcache                                        (hdmi_dmac_0_m_src_axi_arcache),                           //                                                               .arcache
		.hdmi_dmac_0_m_src_axi_arprot                                         (hdmi_dmac_0_m_src_axi_arprot),                            //                                                               .arprot
		.hdmi_dmac_0_m_src_axi_arvalid                                        (hdmi_dmac_0_m_src_axi_arvalid),                           //                                                               .arvalid
		.hdmi_dmac_0_m_src_axi_arready                                        (hdmi_dmac_0_m_src_axi_arready),                           //                                                               .arready
		.hdmi_dmac_0_m_src_axi_rid                                            (hdmi_dmac_0_m_src_axi_rid),                               //                                                               .rid
		.hdmi_dmac_0_m_src_axi_rdata                                          (hdmi_dmac_0_m_src_axi_rdata),                             //                                                               .rdata
		.hdmi_dmac_0_m_src_axi_rresp                                          (hdmi_dmac_0_m_src_axi_rresp),                             //                                                               .rresp
		.hdmi_dmac_0_m_src_axi_rlast                                          (hdmi_dmac_0_m_src_axi_rlast),                             //                                                               .rlast
		.hdmi_dmac_0_m_src_axi_rvalid                                         (hdmi_dmac_0_m_src_axi_rvalid),                            //                                                               .rvalid
		.hdmi_dmac_0_m_src_axi_rready                                         (hdmi_dmac_0_m_src_axi_rready),                            //                                                               .rready
		.sys_hps_h2f_user1_clock_clk                                          (sys_hps_h2f_user1_clock_clk),                             //                                        sys_hps_h2f_user1_clock.clk
		.axi_adc_dma_m_dest_axi_reset_reset_bridge_in_reset_reset             (rst_controller_reset_out_reset),                          //             axi_adc_dma_m_dest_axi_reset_reset_bridge_in_reset.reset
		.sys_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                      // sys_hps_f2h_sdram0_data_translator_reset_reset_bridge_in_reset.reset
		.sys_hps_f2h_sdram0_data_address                                      (mm_interconnect_1_sys_hps_f2h_sdram0_data_address),       //                                        sys_hps_f2h_sdram0_data.address
		.sys_hps_f2h_sdram0_data_write                                        (mm_interconnect_1_sys_hps_f2h_sdram0_data_write),         //                                                               .write
		.sys_hps_f2h_sdram0_data_read                                         (mm_interconnect_1_sys_hps_f2h_sdram0_data_read),          //                                                               .read
		.sys_hps_f2h_sdram0_data_readdata                                     (mm_interconnect_1_sys_hps_f2h_sdram0_data_readdata),      //                                                               .readdata
		.sys_hps_f2h_sdram0_data_writedata                                    (mm_interconnect_1_sys_hps_f2h_sdram0_data_writedata),     //                                                               .writedata
		.sys_hps_f2h_sdram0_data_burstcount                                   (mm_interconnect_1_sys_hps_f2h_sdram0_data_burstcount),    //                                                               .burstcount
		.sys_hps_f2h_sdram0_data_byteenable                                   (mm_interconnect_1_sys_hps_f2h_sdram0_data_byteenable),    //                                                               .byteenable
		.sys_hps_f2h_sdram0_data_readdatavalid                                (mm_interconnect_1_sys_hps_f2h_sdram0_data_readdatavalid), //                                                               .readdatavalid
		.sys_hps_f2h_sdram0_data_waitrequest                                  (mm_interconnect_1_sys_hps_f2h_sdram0_data_waitrequest)    //                                                               .waitrequest
	);

	system_bd_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq), // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq), // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq), // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq), // receiver6.irq
		.sender_irq    (sys_hps_f2h_irq0_irq)      //    sender.irq
	);

	system_bd_irq_mapper_001 irq_mapper_001 (
		.clk        (),                     //       clk.clk
		.reset      (),                     // clk_reset.reset
		.sender_irq (sys_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~sys_rst_reset_n),               // reset_in0.reset
		.clk            (sys_hps_h2f_user1_clock_clk),    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~sys_hps_h2f_reset_reset_n),         // reset_in0.reset
		.clk            (sys_hps_h2f_user1_clock_clk),        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign util_dac_upack_dac_ch_0_data = { util_dac_upack_fifo_rd_data[15:0] };

	assign util_dac_upack_dac_ch_0_data_valid = { util_dac_upack_fifo_rd_valid[0] };

	assign util_dac_upack_dac_ch_1_data = { util_dac_upack_fifo_rd_data[31:16] };

	assign util_dac_upack_dac_ch_1_data_valid = { util_dac_upack_fifo_rd_valid[0] };

	assign util_dac_upack_dac_ch_2_data = { util_dac_upack_fifo_rd_data[47:32] };

	assign util_dac_upack_dac_ch_2_data_valid = { util_dac_upack_fifo_rd_valid[0] };

	assign util_dac_upack_dac_ch_3_data = { util_dac_upack_fifo_rd_data[63:48] };

	assign util_dac_upack_dac_ch_3_data_valid = { util_dac_upack_fifo_rd_valid[0] };

endmodule
