// ghrd_hps_system.v

// Generated using ACDS version 23.2.1 194

`timescale 1 ps / 1 ps
module ghrd_hps_system (
		output wire        emac0_mdio_mac_mdc,          //           emac0_mdio.mac_mdc
		input  wire        emac0_mdio_mac_mdi,          //                     .mac_mdi
		output wire        emac0_mdio_mac_mdo,          //                     .mac_mdo
		output wire        emac0_mdio_mac_mdoe,         //                     .mac_mdoe
		output wire        emac0_app_rst_reset_n,       //        emac0_app_rst.reset_n
		output wire        emac0_mac_tx_clk_o,          //                emac0.mac_tx_clk_o
		input  wire        emac0_mac_tx_clk_i,          //                     .mac_tx_clk_i
		input  wire        emac0_mac_rx_clk,            //                     .mac_rx_clk
		output wire        emac0_mac_rst_tx_n,          //                     .mac_rst_tx_n
		output wire        emac0_mac_rst_rx_n,          //                     .mac_rst_rx_n
		output wire        emac0_mac_txen,              //                     .mac_txen
		output wire        emac0_mac_txer,              //                     .mac_txer
		input  wire        emac0_mac_rxdv,              //                     .mac_rxdv
		input  wire        emac0_mac_rxer,              //                     .mac_rxer
		input  wire [7:0]  emac0_mac_rxd,               //                     .mac_rxd
		input  wire        emac0_mac_col,               //                     .mac_col
		input  wire        emac0_mac_crs,               //                     .mac_crs
		output wire [2:0]  emac0_mac_speed,             //                     .mac_speed
		output wire [7:0]  emac0_mac_txd_o,             //                     .mac_txd_o
		output wire        emac2_app_rst_reset_n,       //        emac2_app_rst.reset_n
		input  wire        spim0_miso_i,                //                spim0.miso_i
		output wire        spim0_mosi_o,                //                     .mosi_o
		output wire        spim0_mosi_oe,               //                     .mosi_oe
		input  wire        spim0_ss_in_n,               //                     .ss_in_n
		output wire        spim0_ss0_n_o,               //                     .ss0_n_o
		output wire        spim0_ss1_n_o,               //                     .ss1_n_o
		output wire        spim0_ss2_n_o,               //                     .ss2_n_o
		output wire        spim0_ss3_n_o,               //                     .ss3_n_o
		output wire        spim0_sclk_out_clk,          //       spim0_sclk_out.clk
		input  wire        i2c1_scl_i_clk,              //           i2c1_scl_i.clk
		output wire        i2c1_scl_oe_clk,             //          i2c1_scl_oe.clk
		input  wire        i2c1_sda_i,                  //                 i2c1.sda_i
		output wire        i2c1_sda_oe,                 //                     .sda_oe
		input  wire        hps_io_hps_osc_clk,          //               hps_io.hps_osc_clk
		inout  wire        hps_io_sdmmc_data0,          //                     .sdmmc_data0
		inout  wire        hps_io_sdmmc_data1,          //                     .sdmmc_data1
		output wire        hps_io_sdmmc_cclk,           //                     .sdmmc_cclk
		inout  wire        hps_io_sdmmc_data2,          //                     .sdmmc_data2
		inout  wire        hps_io_sdmmc_data3,          //                     .sdmmc_data3
		inout  wire        hps_io_sdmmc_cmd,            //                     .sdmmc_cmd
		input  wire        hps_io_usb1_clk,             //                     .usb1_clk
		output wire        hps_io_usb1_stp,             //                     .usb1_stp
		input  wire        hps_io_usb1_dir,             //                     .usb1_dir
		inout  wire        hps_io_usb1_data0,           //                     .usb1_data0
		inout  wire        hps_io_usb1_data1,           //                     .usb1_data1
		input  wire        hps_io_usb1_nxr,             //                     .usb1_nxr
		inout  wire        hps_io_usb1_data2,           //                     .usb1_data2
		inout  wire        hps_io_usb1_data3,           //                     .usb1_data3
		inout  wire        hps_io_usb1_data4,           //                     .usb1_data4
		inout  wire        hps_io_usb1_data5,           //                     .usb1_data5
		inout  wire        hps_io_usb1_data6,           //                     .usb1_data6
		inout  wire        hps_io_usb1_data7,           //                     .usb1_data7
		output wire        hps_io_emac2_tx_clk,         //                     .emac2_tx_clk
		output wire        hps_io_emac2_tx_ctl,         //                     .emac2_tx_ctl
		input  wire        hps_io_emac2_rx_clk,         //                     .emac2_rx_clk
		input  wire        hps_io_emac2_rx_ctl,         //                     .emac2_rx_ctl
		output wire        hps_io_emac2_txd0,           //                     .emac2_txd0
		output wire        hps_io_emac2_txd1,           //                     .emac2_txd1
		input  wire        hps_io_emac2_rxd0,           //                     .emac2_rxd0
		input  wire        hps_io_emac2_rxd1,           //                     .emac2_rxd1
		output wire        hps_io_emac2_txd2,           //                     .emac2_txd2
		output wire        hps_io_emac2_txd3,           //                     .emac2_txd3
		input  wire        hps_io_emac2_rxd2,           //                     .emac2_rxd2
		input  wire        hps_io_emac2_rxd3,           //                     .emac2_rxd3
		inout  wire        hps_io_mdio2_mdio,           //                     .mdio2_mdio
		output wire        hps_io_mdio2_mdc,            //                     .mdio2_mdc
		output wire        hps_io_uart0_tx,             //                     .uart0_tx
		input  wire        hps_io_uart0_rx,             //                     .uart0_rx
		inout  wire        hps_io_i2c0_sda,             //                     .i2c0_sda
		inout  wire        hps_io_i2c0_scl,             //                     .i2c0_scl
		inout  wire        hps_io_gpio6,                //                     .gpio6
		inout  wire        hps_io_gpio7,                //                     .gpio7
		inout  wire        hps_io_gpio8,                //                     .gpio8
		inout  wire        hps_io_gpio9,                //                     .gpio9
		inout  wire        hps_io_gpio10,               //                     .gpio10
		inout  wire        hps_io_gpio11,               //                     .gpio11
		inout  wire        hps_io_gpio28,               //                     .gpio28
		inout  wire        hps_io_gpio34,               //                     .gpio34
		inout  wire        hps_io_gpio35,               //                     .gpio35
		input  wire        usb31_io_vbus_det,           //             usb31_io.vbus_det
		input  wire        usb31_io_flt_bar,            //                     .flt_bar
		output wire [1:0]  usb31_io_usb_ctrl,           //                     .usb_ctrl
		input  wire        usb31_io_usb31_id,           //                     .usb31_id
		input  wire        bank3a_lpddr4_refclk_clk,    // bank3a_lpddr4_refclk.clk
		output wire        bank3a_lpddr4_mem_ck_t,      //        bank3a_lpddr4.mem_ck_t
		output wire        bank3a_lpddr4_mem_ck_c,      //                     .mem_ck_c
		output wire        bank3a_lpddr4_mem_cke,       //                     .mem_cke
		output wire        bank3a_lpddr4_mem_reset_n,   //                     .mem_reset_n
		output wire        bank3a_lpddr4_mem_cs,        //                     .mem_cs
		output wire [5:0]  bank3a_lpddr4_mem_ca,        //                     .mem_ca
		inout  wire [31:0] bank3a_lpddr4_mem_dq,        //                     .mem_dq
		inout  wire [3:0]  bank3a_lpddr4_mem_dqs_t,     //                     .mem_dqs_t
		inout  wire [3:0]  bank3a_lpddr4_mem_dqs_c,     //                     .mem_dqs_c
		inout  wire [3:0]  bank3a_lpddr4_mem_dmi,       //                     .mem_dmi
		input  wire        bank3a_lpddr4_oct_oct_rzqin, //    bank3a_lpddr4_oct.oct_rzqin
		input  wire        sys_reset_reset,             //            sys_reset.reset
		input  wire [1:0]  dipsw_export,                //                dipsw.export
		input  wire [1:0]  pb_export,                   //                   pb.export
		output wire [2:0]  rgb_led0_export,             //             rgb_led0.export
		output wire [2:0]  rgb_led1_export,             //             rgb_led1.export
		output wire [2:0]  rgb_led2_export,             //             rgb_led2.export
		output wire [2:0]  rgb_led3_export,             //             rgb_led3.export
		output wire        hdmi_h_clk,                  //                 hdmi.h_clk
		output wire        hdmi_h16_hsync,              //                     .h16_hsync
		output wire        hdmi_h16_vsync,              //                     .h16_vsync
		output wire        hdmi_h16_data_e,             //                     .h16_data_e
		output wire [15:0] hdmi_h16_data,               //                     .h16_data
		output wire [15:0] hdmi_h16_es_data,            //                     .h16_es_data
		output wire        hdmi_h24_hsync,              //                     .h24_hsync
		output wire        hdmi_h24_vsync,              //                     .h24_vsync
		output wire        hdmi_h24_data_e,             //                     .h24_data_e
		output wire [23:0] hdmi_h24_data,               //                     .h24_data
		output wire        hdmi_h36_hsync,              //                     .h36_hsync
		output wire        hdmi_h36_vsync,              //                     .h36_vsync
		output wire        hdmi_h36_data_e,             //                     .h36_data_e
		output wire [35:0] hdmi_h36_data,               //                     .h36_data
		input  wire        hdmi_pll_refclk_clk          //      hdmi_pll_refclk.clk
	);

	wire          agilex_5_soc_h2f_user0_clk_clk;                                           // agilex_5_soc:h2f_user0_clk_clk -> [agilex_5_soc:emac_ptp_clk_clk, agilex_5_soc:emac_timestamp_clk_clk, mm_interconnect_1:agilex_5_soc_h2f_user0_clk_clk, onchip_sram:clk, rst_controller_003:clk, rst_controller_005:clk]
	wire          agilex_5_soc_h2f_user1_clk_clk;                                           // agilex_5_soc:h2f_user1_clk_clk -> [agilex_5_soc:f2sdram_axi_clock_clk, agilex_5_soc:fpga2hps_clock_clk, agilex_5_soc:hps2fpga_axi_clock_clk, agilex_5_soc:lwhps2fpga_axi_clock_clk, bank3a_emif_master:clk_clk, emif_bank3a:s0_axil_clk, emif_bank3a:usr_async_clk_0, f2sdram_only_master:clk_clk, fpga_only_master:clk_clk, mm_interconnect_0:agilex_5_soc_h2f_user1_clk_clk, mm_interconnect_1:agilex_5_soc_h2f_user1_clk_clk, mm_interconnect_2:agilex_5_soc_h2f_user1_clk_clk, mm_interconnect_3:agilex_5_soc_h2f_user1_clk_clk, peripheral_sys_0:clk_clk, reset_in:clk, rst_controller_001:clk, rst_controller_004:clk, rst_controller_006:clk, rst_controller_007:clk, rst_controller_008:clk, video_sys_0:clk_clk]
	wire          reset_in_out_reset_reset;                                                 // reset_in:out_reset -> [agilex_5_soc:f2sdram_axi_reset_reset_n, agilex_5_soc:fpga2hps_reset_reset_n, agilex_5_soc:hps2fpga_axi_reset_reset_n, agilex_5_soc:lwhps2fpga_axi_reset_reset_n, bank3a_emif_master:clk_reset_reset, f2sdram_only_master:clk_reset_reset, peripheral_sys_0:reset_reset, rst_controller_002:reset_in1, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0, rst_controller_006:reset_in1, video_sys_0:reset_reset]
	wire    [1:0] video_sys_0_hdmi_dmac_master_awburst;                                     // video_sys_0:hdmi_dmac_master_awburst -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awburst
	wire    [3:0] video_sys_0_hdmi_dmac_master_arlen;                                       // video_sys_0:hdmi_dmac_master_arlen -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arlen
	wire    [7:0] video_sys_0_hdmi_dmac_master_wstrb;                                       // video_sys_0:hdmi_dmac_master_wstrb -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_wstrb
	wire          video_sys_0_hdmi_dmac_master_wready;                                      // mm_interconnect_0:video_sys_0_hdmi_dmac_master_wready -> video_sys_0:hdmi_dmac_master_wready
	wire          video_sys_0_hdmi_dmac_master_rid;                                         // mm_interconnect_0:video_sys_0_hdmi_dmac_master_rid -> video_sys_0:hdmi_dmac_master_rid
	wire          video_sys_0_hdmi_dmac_master_rready;                                      // video_sys_0:hdmi_dmac_master_rready -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_rready
	wire    [3:0] video_sys_0_hdmi_dmac_master_awlen;                                       // video_sys_0:hdmi_dmac_master_awlen -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awlen
	wire          video_sys_0_hdmi_dmac_master_wid;                                         // video_sys_0:hdmi_dmac_master_wid -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_wid
	wire    [3:0] video_sys_0_hdmi_dmac_master_arcache;                                     // video_sys_0:hdmi_dmac_master_arcache -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arcache
	wire          video_sys_0_hdmi_dmac_master_wvalid;                                      // video_sys_0:hdmi_dmac_master_wvalid -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_wvalid
	wire   [31:0] video_sys_0_hdmi_dmac_master_araddr;                                      // video_sys_0:hdmi_dmac_master_araddr -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_araddr
	wire    [2:0] video_sys_0_hdmi_dmac_master_arprot;                                      // video_sys_0:hdmi_dmac_master_arprot -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arprot
	wire   [63:0] video_sys_0_hdmi_dmac_master_wdata;                                       // video_sys_0:hdmi_dmac_master_wdata -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_wdata
	wire          video_sys_0_hdmi_dmac_master_arvalid;                                     // video_sys_0:hdmi_dmac_master_arvalid -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arvalid
	wire    [2:0] video_sys_0_hdmi_dmac_master_awprot;                                      // video_sys_0:hdmi_dmac_master_awprot -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awprot
	wire    [3:0] video_sys_0_hdmi_dmac_master_awcache;                                     // video_sys_0:hdmi_dmac_master_awcache -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awcache
	wire          video_sys_0_hdmi_dmac_master_arid;                                        // video_sys_0:hdmi_dmac_master_arid -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arid
	wire    [1:0] video_sys_0_hdmi_dmac_master_arlock;                                      // video_sys_0:hdmi_dmac_master_arlock -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arlock
	wire    [1:0] video_sys_0_hdmi_dmac_master_awlock;                                      // video_sys_0:hdmi_dmac_master_awlock -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awlock
	wire   [31:0] video_sys_0_hdmi_dmac_master_awaddr;                                      // video_sys_0:hdmi_dmac_master_awaddr -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awaddr
	wire    [1:0] video_sys_0_hdmi_dmac_master_bresp;                                       // mm_interconnect_0:video_sys_0_hdmi_dmac_master_bresp -> video_sys_0:hdmi_dmac_master_bresp
	wire          video_sys_0_hdmi_dmac_master_arready;                                     // mm_interconnect_0:video_sys_0_hdmi_dmac_master_arready -> video_sys_0:hdmi_dmac_master_arready
	wire   [63:0] video_sys_0_hdmi_dmac_master_rdata;                                       // mm_interconnect_0:video_sys_0_hdmi_dmac_master_rdata -> video_sys_0:hdmi_dmac_master_rdata
	wire          video_sys_0_hdmi_dmac_master_awready;                                     // mm_interconnect_0:video_sys_0_hdmi_dmac_master_awready -> video_sys_0:hdmi_dmac_master_awready
	wire    [1:0] video_sys_0_hdmi_dmac_master_arburst;                                     // video_sys_0:hdmi_dmac_master_arburst -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arburst
	wire    [2:0] video_sys_0_hdmi_dmac_master_arsize;                                      // video_sys_0:hdmi_dmac_master_arsize -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_arsize
	wire          video_sys_0_hdmi_dmac_master_bready;                                      // video_sys_0:hdmi_dmac_master_bready -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_bready
	wire          video_sys_0_hdmi_dmac_master_rlast;                                       // mm_interconnect_0:video_sys_0_hdmi_dmac_master_rlast -> video_sys_0:hdmi_dmac_master_rlast
	wire          video_sys_0_hdmi_dmac_master_wlast;                                       // video_sys_0:hdmi_dmac_master_wlast -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_wlast
	wire    [1:0] video_sys_0_hdmi_dmac_master_rresp;                                       // mm_interconnect_0:video_sys_0_hdmi_dmac_master_rresp -> video_sys_0:hdmi_dmac_master_rresp
	wire          video_sys_0_hdmi_dmac_master_awid;                                        // video_sys_0:hdmi_dmac_master_awid -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awid
	wire          video_sys_0_hdmi_dmac_master_bid;                                         // mm_interconnect_0:video_sys_0_hdmi_dmac_master_bid -> video_sys_0:hdmi_dmac_master_bid
	wire          video_sys_0_hdmi_dmac_master_bvalid;                                      // mm_interconnect_0:video_sys_0_hdmi_dmac_master_bvalid -> video_sys_0:hdmi_dmac_master_bvalid
	wire          video_sys_0_hdmi_dmac_master_awvalid;                                     // video_sys_0:hdmi_dmac_master_awvalid -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awvalid
	wire          video_sys_0_hdmi_dmac_master_rvalid;                                      // mm_interconnect_0:video_sys_0_hdmi_dmac_master_rvalid -> video_sys_0:hdmi_dmac_master_rvalid
	wire    [2:0] video_sys_0_hdmi_dmac_master_awsize;                                      // video_sys_0:hdmi_dmac_master_awsize -> mm_interconnect_0:video_sys_0_hdmi_dmac_master_awsize
	wire   [31:0] f2sdram_only_master_master_readdata;                                      // mm_interconnect_0:f2sdram_only_master_master_readdata -> f2sdram_only_master:master_readdata
	wire          f2sdram_only_master_master_waitrequest;                                   // mm_interconnect_0:f2sdram_only_master_master_waitrequest -> f2sdram_only_master:master_waitrequest
	wire   [31:0] f2sdram_only_master_master_address;                                       // f2sdram_only_master:master_address -> mm_interconnect_0:f2sdram_only_master_master_address
	wire          f2sdram_only_master_master_read;                                          // f2sdram_only_master:master_read -> mm_interconnect_0:f2sdram_only_master_master_read
	wire    [3:0] f2sdram_only_master_master_byteenable;                                    // f2sdram_only_master:master_byteenable -> mm_interconnect_0:f2sdram_only_master_master_byteenable
	wire          f2sdram_only_master_master_readdatavalid;                                 // mm_interconnect_0:f2sdram_only_master_master_readdatavalid -> f2sdram_only_master:master_readdatavalid
	wire          f2sdram_only_master_master_write;                                         // f2sdram_only_master:master_write -> mm_interconnect_0:f2sdram_only_master_master_write
	wire   [31:0] f2sdram_only_master_master_writedata;                                     // f2sdram_only_master:master_writedata -> mm_interconnect_0:f2sdram_only_master_master_writedata
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_ruser;                             // agilex_5_soc:f2sdram_ruser -> mm_interconnect_0:agilex_5_soc_f2sdram_ruser
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_wuser;                             // mm_interconnect_0:agilex_5_soc_f2sdram_wuser -> agilex_5_soc:f2sdram_wuser
	wire    [1:0] mm_interconnect_0_agilex_5_soc_f2sdram_awburst;                           // mm_interconnect_0:agilex_5_soc_f2sdram_awburst -> agilex_5_soc:f2sdram_awburst
	wire    [3:0] mm_interconnect_0_agilex_5_soc_f2sdram_arregion;                          // mm_interconnect_0:agilex_5_soc_f2sdram_arregion -> agilex_5_soc:f2sdram_arregion
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_awuser;                            // mm_interconnect_0:agilex_5_soc_f2sdram_awuser -> agilex_5_soc:f2sdram_awuser
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_arlen;                             // mm_interconnect_0:agilex_5_soc_f2sdram_arlen -> agilex_5_soc:f2sdram_arlen
	wire    [3:0] mm_interconnect_0_agilex_5_soc_f2sdram_arqos;                             // mm_interconnect_0:agilex_5_soc_f2sdram_arqos -> agilex_5_soc:f2sdram_arqos
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_wstrb;                             // mm_interconnect_0:agilex_5_soc_f2sdram_wstrb -> agilex_5_soc:f2sdram_wstrb
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_wready;                            // agilex_5_soc:f2sdram_wready -> mm_interconnect_0:agilex_5_soc_f2sdram_wready
	wire    [4:0] mm_interconnect_0_agilex_5_soc_f2sdram_rid;                               // agilex_5_soc:f2sdram_rid -> mm_interconnect_0:agilex_5_soc_f2sdram_rid
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_rready;                            // mm_interconnect_0:agilex_5_soc_f2sdram_rready -> agilex_5_soc:f2sdram_rready
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_awlen;                             // mm_interconnect_0:agilex_5_soc_f2sdram_awlen -> agilex_5_soc:f2sdram_awlen
	wire    [3:0] mm_interconnect_0_agilex_5_soc_f2sdram_awqos;                             // mm_interconnect_0:agilex_5_soc_f2sdram_awqos -> agilex_5_soc:f2sdram_awqos
	wire    [3:0] mm_interconnect_0_agilex_5_soc_f2sdram_arcache;                           // mm_interconnect_0:agilex_5_soc_f2sdram_arcache -> agilex_5_soc:f2sdram_arcache
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_wvalid;                            // mm_interconnect_0:agilex_5_soc_f2sdram_wvalid -> agilex_5_soc:f2sdram_wvalid
	wire   [31:0] mm_interconnect_0_agilex_5_soc_f2sdram_araddr;                            // mm_interconnect_0:agilex_5_soc_f2sdram_araddr -> agilex_5_soc:f2sdram_araddr
	wire    [2:0] mm_interconnect_0_agilex_5_soc_f2sdram_arprot;                            // mm_interconnect_0:agilex_5_soc_f2sdram_arprot -> agilex_5_soc:f2sdram_arprot
	wire    [2:0] mm_interconnect_0_agilex_5_soc_f2sdram_awprot;                            // mm_interconnect_0:agilex_5_soc_f2sdram_awprot -> agilex_5_soc:f2sdram_awprot
	wire   [63:0] mm_interconnect_0_agilex_5_soc_f2sdram_wdata;                             // mm_interconnect_0:agilex_5_soc_f2sdram_wdata -> agilex_5_soc:f2sdram_wdata
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_arvalid;                           // mm_interconnect_0:agilex_5_soc_f2sdram_arvalid -> agilex_5_soc:f2sdram_arvalid
	wire    [3:0] mm_interconnect_0_agilex_5_soc_f2sdram_awcache;                           // mm_interconnect_0:agilex_5_soc_f2sdram_awcache -> agilex_5_soc:f2sdram_awcache
	wire    [4:0] mm_interconnect_0_agilex_5_soc_f2sdram_arid;                              // mm_interconnect_0:agilex_5_soc_f2sdram_arid -> agilex_5_soc:f2sdram_arid
	wire    [0:0] mm_interconnect_0_agilex_5_soc_f2sdram_arlock;                            // mm_interconnect_0:agilex_5_soc_f2sdram_arlock -> agilex_5_soc:f2sdram_arlock
	wire    [0:0] mm_interconnect_0_agilex_5_soc_f2sdram_awlock;                            // mm_interconnect_0:agilex_5_soc_f2sdram_awlock -> agilex_5_soc:f2sdram_awlock
	wire   [31:0] mm_interconnect_0_agilex_5_soc_f2sdram_awaddr;                            // mm_interconnect_0:agilex_5_soc_f2sdram_awaddr -> agilex_5_soc:f2sdram_awaddr
	wire    [1:0] mm_interconnect_0_agilex_5_soc_f2sdram_bresp;                             // agilex_5_soc:f2sdram_bresp -> mm_interconnect_0:agilex_5_soc_f2sdram_bresp
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_arready;                           // agilex_5_soc:f2sdram_arready -> mm_interconnect_0:agilex_5_soc_f2sdram_arready
	wire   [63:0] mm_interconnect_0_agilex_5_soc_f2sdram_rdata;                             // agilex_5_soc:f2sdram_rdata -> mm_interconnect_0:agilex_5_soc_f2sdram_rdata
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_awready;                           // agilex_5_soc:f2sdram_awready -> mm_interconnect_0:agilex_5_soc_f2sdram_awready
	wire    [1:0] mm_interconnect_0_agilex_5_soc_f2sdram_arburst;                           // mm_interconnect_0:agilex_5_soc_f2sdram_arburst -> agilex_5_soc:f2sdram_arburst
	wire    [2:0] mm_interconnect_0_agilex_5_soc_f2sdram_arsize;                            // mm_interconnect_0:agilex_5_soc_f2sdram_arsize -> agilex_5_soc:f2sdram_arsize
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_bready;                            // mm_interconnect_0:agilex_5_soc_f2sdram_bready -> agilex_5_soc:f2sdram_bready
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_rlast;                             // agilex_5_soc:f2sdram_rlast -> mm_interconnect_0:agilex_5_soc_f2sdram_rlast
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_wlast;                             // mm_interconnect_0:agilex_5_soc_f2sdram_wlast -> agilex_5_soc:f2sdram_wlast
	wire    [3:0] mm_interconnect_0_agilex_5_soc_f2sdram_awregion;                          // mm_interconnect_0:agilex_5_soc_f2sdram_awregion -> agilex_5_soc:f2sdram_awregion
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_buser;                             // agilex_5_soc:f2sdram_buser -> mm_interconnect_0:agilex_5_soc_f2sdram_buser
	wire    [1:0] mm_interconnect_0_agilex_5_soc_f2sdram_rresp;                             // agilex_5_soc:f2sdram_rresp -> mm_interconnect_0:agilex_5_soc_f2sdram_rresp
	wire    [4:0] mm_interconnect_0_agilex_5_soc_f2sdram_awid;                              // mm_interconnect_0:agilex_5_soc_f2sdram_awid -> agilex_5_soc:f2sdram_awid
	wire    [4:0] mm_interconnect_0_agilex_5_soc_f2sdram_bid;                               // agilex_5_soc:f2sdram_bid -> mm_interconnect_0:agilex_5_soc_f2sdram_bid
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_bvalid;                            // agilex_5_soc:f2sdram_bvalid -> mm_interconnect_0:agilex_5_soc_f2sdram_bvalid
	wire    [2:0] mm_interconnect_0_agilex_5_soc_f2sdram_awsize;                            // mm_interconnect_0:agilex_5_soc_f2sdram_awsize -> agilex_5_soc:f2sdram_awsize
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_awvalid;                           // mm_interconnect_0:agilex_5_soc_f2sdram_awvalid -> agilex_5_soc:f2sdram_awvalid
	wire    [7:0] mm_interconnect_0_agilex_5_soc_f2sdram_aruser;                            // mm_interconnect_0:agilex_5_soc_f2sdram_aruser -> agilex_5_soc:f2sdram_aruser
	wire          mm_interconnect_0_agilex_5_soc_f2sdram_rvalid;                            // agilex_5_soc:f2sdram_rvalid -> mm_interconnect_0:agilex_5_soc_f2sdram_rvalid
	wire    [1:0] agilex_5_soc_hps2fpga_awburst;                                            // agilex_5_soc:hps2fpga_awburst -> mm_interconnect_1:agilex_5_soc_hps2fpga_awburst
	wire    [7:0] agilex_5_soc_hps2fpga_arlen;                                              // agilex_5_soc:hps2fpga_arlen -> mm_interconnect_1:agilex_5_soc_hps2fpga_arlen
	wire    [3:0] agilex_5_soc_hps2fpga_wstrb;                                              // agilex_5_soc:hps2fpga_wstrb -> mm_interconnect_1:agilex_5_soc_hps2fpga_wstrb
	wire          agilex_5_soc_hps2fpga_wready;                                             // mm_interconnect_1:agilex_5_soc_hps2fpga_wready -> agilex_5_soc:hps2fpga_wready
	wire    [3:0] agilex_5_soc_hps2fpga_rid;                                                // mm_interconnect_1:agilex_5_soc_hps2fpga_rid -> agilex_5_soc:hps2fpga_rid
	wire          agilex_5_soc_hps2fpga_rready;                                             // agilex_5_soc:hps2fpga_rready -> mm_interconnect_1:agilex_5_soc_hps2fpga_rready
	wire    [7:0] agilex_5_soc_hps2fpga_awlen;                                              // agilex_5_soc:hps2fpga_awlen -> mm_interconnect_1:agilex_5_soc_hps2fpga_awlen
	wire    [3:0] agilex_5_soc_hps2fpga_arcache;                                            // agilex_5_soc:hps2fpga_arcache -> mm_interconnect_1:agilex_5_soc_hps2fpga_arcache
	wire          agilex_5_soc_hps2fpga_wvalid;                                             // agilex_5_soc:hps2fpga_wvalid -> mm_interconnect_1:agilex_5_soc_hps2fpga_wvalid
	wire   [31:0] agilex_5_soc_hps2fpga_araddr;                                             // agilex_5_soc:hps2fpga_araddr -> mm_interconnect_1:agilex_5_soc_hps2fpga_araddr
	wire    [2:0] agilex_5_soc_hps2fpga_arprot;                                             // agilex_5_soc:hps2fpga_arprot -> mm_interconnect_1:agilex_5_soc_hps2fpga_arprot
	wire    [2:0] agilex_5_soc_hps2fpga_awprot;                                             // agilex_5_soc:hps2fpga_awprot -> mm_interconnect_1:agilex_5_soc_hps2fpga_awprot
	wire   [31:0] agilex_5_soc_hps2fpga_wdata;                                              // agilex_5_soc:hps2fpga_wdata -> mm_interconnect_1:agilex_5_soc_hps2fpga_wdata
	wire          agilex_5_soc_hps2fpga_arvalid;                                            // agilex_5_soc:hps2fpga_arvalid -> mm_interconnect_1:agilex_5_soc_hps2fpga_arvalid
	wire    [3:0] agilex_5_soc_hps2fpga_awcache;                                            // agilex_5_soc:hps2fpga_awcache -> mm_interconnect_1:agilex_5_soc_hps2fpga_awcache
	wire    [3:0] agilex_5_soc_hps2fpga_arid;                                               // agilex_5_soc:hps2fpga_arid -> mm_interconnect_1:agilex_5_soc_hps2fpga_arid
	wire          agilex_5_soc_hps2fpga_arlock;                                             // agilex_5_soc:hps2fpga_arlock -> mm_interconnect_1:agilex_5_soc_hps2fpga_arlock
	wire          agilex_5_soc_hps2fpga_awlock;                                             // agilex_5_soc:hps2fpga_awlock -> mm_interconnect_1:agilex_5_soc_hps2fpga_awlock
	wire   [31:0] agilex_5_soc_hps2fpga_awaddr;                                             // agilex_5_soc:hps2fpga_awaddr -> mm_interconnect_1:agilex_5_soc_hps2fpga_awaddr
	wire    [1:0] agilex_5_soc_hps2fpga_bresp;                                              // mm_interconnect_1:agilex_5_soc_hps2fpga_bresp -> agilex_5_soc:hps2fpga_bresp
	wire          agilex_5_soc_hps2fpga_arready;                                            // mm_interconnect_1:agilex_5_soc_hps2fpga_arready -> agilex_5_soc:hps2fpga_arready
	wire   [31:0] agilex_5_soc_hps2fpga_rdata;                                              // mm_interconnect_1:agilex_5_soc_hps2fpga_rdata -> agilex_5_soc:hps2fpga_rdata
	wire          agilex_5_soc_hps2fpga_awready;                                            // mm_interconnect_1:agilex_5_soc_hps2fpga_awready -> agilex_5_soc:hps2fpga_awready
	wire    [1:0] agilex_5_soc_hps2fpga_arburst;                                            // agilex_5_soc:hps2fpga_arburst -> mm_interconnect_1:agilex_5_soc_hps2fpga_arburst
	wire    [2:0] agilex_5_soc_hps2fpga_arsize;                                             // agilex_5_soc:hps2fpga_arsize -> mm_interconnect_1:agilex_5_soc_hps2fpga_arsize
	wire          agilex_5_soc_hps2fpga_bready;                                             // agilex_5_soc:hps2fpga_bready -> mm_interconnect_1:agilex_5_soc_hps2fpga_bready
	wire          agilex_5_soc_hps2fpga_rlast;                                              // mm_interconnect_1:agilex_5_soc_hps2fpga_rlast -> agilex_5_soc:hps2fpga_rlast
	wire          agilex_5_soc_hps2fpga_wlast;                                              // agilex_5_soc:hps2fpga_wlast -> mm_interconnect_1:agilex_5_soc_hps2fpga_wlast
	wire    [1:0] agilex_5_soc_hps2fpga_rresp;                                              // mm_interconnect_1:agilex_5_soc_hps2fpga_rresp -> agilex_5_soc:hps2fpga_rresp
	wire    [3:0] agilex_5_soc_hps2fpga_awid;                                               // agilex_5_soc:hps2fpga_awid -> mm_interconnect_1:agilex_5_soc_hps2fpga_awid
	wire    [3:0] agilex_5_soc_hps2fpga_bid;                                                // mm_interconnect_1:agilex_5_soc_hps2fpga_bid -> agilex_5_soc:hps2fpga_bid
	wire          agilex_5_soc_hps2fpga_bvalid;                                             // mm_interconnect_1:agilex_5_soc_hps2fpga_bvalid -> agilex_5_soc:hps2fpga_bvalid
	wire    [2:0] agilex_5_soc_hps2fpga_awsize;                                             // agilex_5_soc:hps2fpga_awsize -> mm_interconnect_1:agilex_5_soc_hps2fpga_awsize
	wire          agilex_5_soc_hps2fpga_awvalid;                                            // agilex_5_soc:hps2fpga_awvalid -> mm_interconnect_1:agilex_5_soc_hps2fpga_awvalid
	wire          agilex_5_soc_hps2fpga_rvalid;                                             // mm_interconnect_1:agilex_5_soc_hps2fpga_rvalid -> agilex_5_soc:hps2fpga_rvalid
	wire   [31:0] fpga_only_master_master_readdata;                                         // mm_interconnect_1:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	wire          fpga_only_master_master_waitrequest;                                      // mm_interconnect_1:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	wire   [31:0] fpga_only_master_master_address;                                          // fpga_only_master:master_address -> mm_interconnect_1:fpga_only_master_master_address
	wire          fpga_only_master_master_read;                                             // fpga_only_master:master_read -> mm_interconnect_1:fpga_only_master_master_read
	wire    [3:0] fpga_only_master_master_byteenable;                                       // fpga_only_master:master_byteenable -> mm_interconnect_1:fpga_only_master_master_byteenable
	wire          fpga_only_master_master_readdatavalid;                                    // mm_interconnect_1:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	wire          fpga_only_master_master_write;                                            // fpga_only_master:master_write -> mm_interconnect_1:fpga_only_master_master_write
	wire   [31:0] fpga_only_master_master_writedata;                                        // fpga_only_master:master_writedata -> mm_interconnect_1:fpga_only_master_master_writedata
	wire    [1:0] mm_interconnect_1_onchip_sram_axi_s1_awburst;                             // mm_interconnect_1:onchip_sram_axi_s1_awburst -> onchip_sram:s1_awburst
	wire    [7:0] mm_interconnect_1_onchip_sram_axi_s1_arlen;                               // mm_interconnect_1:onchip_sram_axi_s1_arlen -> onchip_sram:s1_arlen
	wire    [7:0] mm_interconnect_1_onchip_sram_axi_s1_wstrb;                               // mm_interconnect_1:onchip_sram_axi_s1_wstrb -> onchip_sram:s1_wstrb
	wire          mm_interconnect_1_onchip_sram_axi_s1_wready;                              // onchip_sram:s1_wready -> mm_interconnect_1:onchip_sram_axi_s1_wready
	wire    [6:0] mm_interconnect_1_onchip_sram_axi_s1_rid;                                 // onchip_sram:s1_rid -> mm_interconnect_1:onchip_sram_axi_s1_rid
	wire          mm_interconnect_1_onchip_sram_axi_s1_rready;                              // mm_interconnect_1:onchip_sram_axi_s1_rready -> onchip_sram:s1_rready
	wire    [7:0] mm_interconnect_1_onchip_sram_axi_s1_awlen;                               // mm_interconnect_1:onchip_sram_axi_s1_awlen -> onchip_sram:s1_awlen
	wire          mm_interconnect_1_onchip_sram_axi_s1_wvalid;                              // mm_interconnect_1:onchip_sram_axi_s1_wvalid -> onchip_sram:s1_wvalid
	wire   [14:0] mm_interconnect_1_onchip_sram_axi_s1_araddr;                              // mm_interconnect_1:onchip_sram_axi_s1_araddr -> onchip_sram:s1_araddr
	wire   [63:0] mm_interconnect_1_onchip_sram_axi_s1_wdata;                               // mm_interconnect_1:onchip_sram_axi_s1_wdata -> onchip_sram:s1_wdata
	wire          mm_interconnect_1_onchip_sram_axi_s1_arvalid;                             // mm_interconnect_1:onchip_sram_axi_s1_arvalid -> onchip_sram:s1_arvalid
	wire    [6:0] mm_interconnect_1_onchip_sram_axi_s1_arid;                                // mm_interconnect_1:onchip_sram_axi_s1_arid -> onchip_sram:s1_arid
	wire   [14:0] mm_interconnect_1_onchip_sram_axi_s1_awaddr;                              // mm_interconnect_1:onchip_sram_axi_s1_awaddr -> onchip_sram:s1_awaddr
	wire    [1:0] mm_interconnect_1_onchip_sram_axi_s1_bresp;                               // onchip_sram:s1_bresp -> mm_interconnect_1:onchip_sram_axi_s1_bresp
	wire          mm_interconnect_1_onchip_sram_axi_s1_arready;                             // onchip_sram:s1_arready -> mm_interconnect_1:onchip_sram_axi_s1_arready
	wire   [63:0] mm_interconnect_1_onchip_sram_axi_s1_rdata;                               // onchip_sram:s1_rdata -> mm_interconnect_1:onchip_sram_axi_s1_rdata
	wire          mm_interconnect_1_onchip_sram_axi_s1_awready;                             // onchip_sram:s1_awready -> mm_interconnect_1:onchip_sram_axi_s1_awready
	wire    [1:0] mm_interconnect_1_onchip_sram_axi_s1_arburst;                             // mm_interconnect_1:onchip_sram_axi_s1_arburst -> onchip_sram:s1_arburst
	wire    [2:0] mm_interconnect_1_onchip_sram_axi_s1_arsize;                              // mm_interconnect_1:onchip_sram_axi_s1_arsize -> onchip_sram:s1_arsize
	wire          mm_interconnect_1_onchip_sram_axi_s1_bready;                              // mm_interconnect_1:onchip_sram_axi_s1_bready -> onchip_sram:s1_bready
	wire          mm_interconnect_1_onchip_sram_axi_s1_rlast;                               // onchip_sram:s1_rlast -> mm_interconnect_1:onchip_sram_axi_s1_rlast
	wire          mm_interconnect_1_onchip_sram_axi_s1_wlast;                               // mm_interconnect_1:onchip_sram_axi_s1_wlast -> onchip_sram:s1_wlast
	wire    [1:0] mm_interconnect_1_onchip_sram_axi_s1_rresp;                               // onchip_sram:s1_rresp -> mm_interconnect_1:onchip_sram_axi_s1_rresp
	wire    [6:0] mm_interconnect_1_onchip_sram_axi_s1_awid;                                // mm_interconnect_1:onchip_sram_axi_s1_awid -> onchip_sram:s1_awid
	wire    [6:0] mm_interconnect_1_onchip_sram_axi_s1_bid;                                 // onchip_sram:s1_bid -> mm_interconnect_1:onchip_sram_axi_s1_bid
	wire          mm_interconnect_1_onchip_sram_axi_s1_bvalid;                              // onchip_sram:s1_bvalid -> mm_interconnect_1:onchip_sram_axi_s1_bvalid
	wire    [2:0] mm_interconnect_1_onchip_sram_axi_s1_awsize;                              // mm_interconnect_1:onchip_sram_axi_s1_awsize -> onchip_sram:s1_awsize
	wire          mm_interconnect_1_onchip_sram_axi_s1_awvalid;                             // mm_interconnect_1:onchip_sram_axi_s1_awvalid -> onchip_sram:s1_awvalid
	wire          mm_interconnect_1_onchip_sram_axi_s1_rvalid;                              // onchip_sram:s1_rvalid -> mm_interconnect_1:onchip_sram_axi_s1_rvalid
	wire   [31:0] mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_readdata;      // peripheral_sys_0:mm_peripheral_bridge_s0_readdata -> mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_readdata
	wire          mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_waitrequest;   // peripheral_sys_0:mm_peripheral_bridge_s0_waitrequest -> mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_waitrequest
	wire          mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_debugaccess;   // mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_debugaccess -> peripheral_sys_0:mm_peripheral_bridge_s0_debugaccess
	wire   [23:0] mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_address;       // mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_address -> peripheral_sys_0:mm_peripheral_bridge_s0_address
	wire          mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_read;          // mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_read -> peripheral_sys_0:mm_peripheral_bridge_s0_read
	wire    [3:0] mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_byteenable;    // mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_byteenable -> peripheral_sys_0:mm_peripheral_bridge_s0_byteenable
	wire          mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_readdatavalid; // peripheral_sys_0:mm_peripheral_bridge_s0_readdatavalid -> mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_readdatavalid
	wire          mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_write;         // mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_write -> peripheral_sys_0:mm_peripheral_bridge_s0_write
	wire   [31:0] mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_writedata;     // mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_writedata -> peripheral_sys_0:mm_peripheral_bridge_s0_writedata
	wire    [0:0] mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_burstcount;    // mm_interconnect_1:peripheral_sys_0_mm_peripheral_bridge_s0_burstcount -> peripheral_sys_0:mm_peripheral_bridge_s0_burstcount
	wire    [1:0] agilex_5_soc_lwhps2fpga_awburst;                                          // agilex_5_soc:lwhps2fpga_awburst -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awburst
	wire    [7:0] agilex_5_soc_lwhps2fpga_arlen;                                            // agilex_5_soc:lwhps2fpga_arlen -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arlen
	wire    [3:0] agilex_5_soc_lwhps2fpga_wstrb;                                            // agilex_5_soc:lwhps2fpga_wstrb -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_wstrb
	wire          agilex_5_soc_lwhps2fpga_wready;                                           // mm_interconnect_2:agilex_5_soc_lwhps2fpga_wready -> agilex_5_soc:lwhps2fpga_wready
	wire    [3:0] agilex_5_soc_lwhps2fpga_rid;                                              // mm_interconnect_2:agilex_5_soc_lwhps2fpga_rid -> agilex_5_soc:lwhps2fpga_rid
	wire          agilex_5_soc_lwhps2fpga_rready;                                           // agilex_5_soc:lwhps2fpga_rready -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_rready
	wire    [7:0] agilex_5_soc_lwhps2fpga_awlen;                                            // agilex_5_soc:lwhps2fpga_awlen -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awlen
	wire    [3:0] agilex_5_soc_lwhps2fpga_arcache;                                          // agilex_5_soc:lwhps2fpga_arcache -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arcache
	wire          agilex_5_soc_lwhps2fpga_wvalid;                                           // agilex_5_soc:lwhps2fpga_wvalid -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_wvalid
	wire   [28:0] agilex_5_soc_lwhps2fpga_araddr;                                           // agilex_5_soc:lwhps2fpga_araddr -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_araddr
	wire    [2:0] agilex_5_soc_lwhps2fpga_arprot;                                           // agilex_5_soc:lwhps2fpga_arprot -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arprot
	wire    [2:0] agilex_5_soc_lwhps2fpga_awprot;                                           // agilex_5_soc:lwhps2fpga_awprot -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awprot
	wire   [31:0] agilex_5_soc_lwhps2fpga_wdata;                                            // agilex_5_soc:lwhps2fpga_wdata -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_wdata
	wire          agilex_5_soc_lwhps2fpga_arvalid;                                          // agilex_5_soc:lwhps2fpga_arvalid -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arvalid
	wire    [3:0] agilex_5_soc_lwhps2fpga_awcache;                                          // agilex_5_soc:lwhps2fpga_awcache -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awcache
	wire    [3:0] agilex_5_soc_lwhps2fpga_arid;                                             // agilex_5_soc:lwhps2fpga_arid -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arid
	wire          agilex_5_soc_lwhps2fpga_arlock;                                           // agilex_5_soc:lwhps2fpga_arlock -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arlock
	wire          agilex_5_soc_lwhps2fpga_awlock;                                           // agilex_5_soc:lwhps2fpga_awlock -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awlock
	wire   [28:0] agilex_5_soc_lwhps2fpga_awaddr;                                           // agilex_5_soc:lwhps2fpga_awaddr -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awaddr
	wire    [1:0] agilex_5_soc_lwhps2fpga_bresp;                                            // mm_interconnect_2:agilex_5_soc_lwhps2fpga_bresp -> agilex_5_soc:lwhps2fpga_bresp
	wire          agilex_5_soc_lwhps2fpga_arready;                                          // mm_interconnect_2:agilex_5_soc_lwhps2fpga_arready -> agilex_5_soc:lwhps2fpga_arready
	wire   [31:0] agilex_5_soc_lwhps2fpga_rdata;                                            // mm_interconnect_2:agilex_5_soc_lwhps2fpga_rdata -> agilex_5_soc:lwhps2fpga_rdata
	wire          agilex_5_soc_lwhps2fpga_awready;                                          // mm_interconnect_2:agilex_5_soc_lwhps2fpga_awready -> agilex_5_soc:lwhps2fpga_awready
	wire    [1:0] agilex_5_soc_lwhps2fpga_arburst;                                          // agilex_5_soc:lwhps2fpga_arburst -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arburst
	wire    [2:0] agilex_5_soc_lwhps2fpga_arsize;                                           // agilex_5_soc:lwhps2fpga_arsize -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_arsize
	wire          agilex_5_soc_lwhps2fpga_bready;                                           // agilex_5_soc:lwhps2fpga_bready -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_bready
	wire          agilex_5_soc_lwhps2fpga_rlast;                                            // mm_interconnect_2:agilex_5_soc_lwhps2fpga_rlast -> agilex_5_soc:lwhps2fpga_rlast
	wire          agilex_5_soc_lwhps2fpga_wlast;                                            // agilex_5_soc:lwhps2fpga_wlast -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_wlast
	wire    [1:0] agilex_5_soc_lwhps2fpga_rresp;                                            // mm_interconnect_2:agilex_5_soc_lwhps2fpga_rresp -> agilex_5_soc:lwhps2fpga_rresp
	wire    [3:0] agilex_5_soc_lwhps2fpga_awid;                                             // agilex_5_soc:lwhps2fpga_awid -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awid
	wire    [3:0] agilex_5_soc_lwhps2fpga_bid;                                              // mm_interconnect_2:agilex_5_soc_lwhps2fpga_bid -> agilex_5_soc:lwhps2fpga_bid
	wire          agilex_5_soc_lwhps2fpga_bvalid;                                           // mm_interconnect_2:agilex_5_soc_lwhps2fpga_bvalid -> agilex_5_soc:lwhps2fpga_bvalid
	wire    [2:0] agilex_5_soc_lwhps2fpga_awsize;                                           // agilex_5_soc:lwhps2fpga_awsize -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awsize
	wire          agilex_5_soc_lwhps2fpga_awvalid;                                          // agilex_5_soc:lwhps2fpga_awvalid -> mm_interconnect_2:agilex_5_soc_lwhps2fpga_awvalid
	wire          agilex_5_soc_lwhps2fpga_rvalid;                                           // mm_interconnect_2:agilex_5_soc_lwhps2fpga_rvalid -> agilex_5_soc:lwhps2fpga_rvalid
	wire   [31:0] mm_interconnect_2_video_sys_0_mm_video_bridge_s0_readdata;                // video_sys_0:mm_video_bridge_s0_readdata -> mm_interconnect_2:video_sys_0_mm_video_bridge_s0_readdata
	wire          mm_interconnect_2_video_sys_0_mm_video_bridge_s0_waitrequest;             // video_sys_0:mm_video_bridge_s0_waitrequest -> mm_interconnect_2:video_sys_0_mm_video_bridge_s0_waitrequest
	wire          mm_interconnect_2_video_sys_0_mm_video_bridge_s0_debugaccess;             // mm_interconnect_2:video_sys_0_mm_video_bridge_s0_debugaccess -> video_sys_0:mm_video_bridge_s0_debugaccess
	wire   [23:0] mm_interconnect_2_video_sys_0_mm_video_bridge_s0_address;                 // mm_interconnect_2:video_sys_0_mm_video_bridge_s0_address -> video_sys_0:mm_video_bridge_s0_address
	wire          mm_interconnect_2_video_sys_0_mm_video_bridge_s0_read;                    // mm_interconnect_2:video_sys_0_mm_video_bridge_s0_read -> video_sys_0:mm_video_bridge_s0_read
	wire    [3:0] mm_interconnect_2_video_sys_0_mm_video_bridge_s0_byteenable;              // mm_interconnect_2:video_sys_0_mm_video_bridge_s0_byteenable -> video_sys_0:mm_video_bridge_s0_byteenable
	wire          mm_interconnect_2_video_sys_0_mm_video_bridge_s0_readdatavalid;           // video_sys_0:mm_video_bridge_s0_readdatavalid -> mm_interconnect_2:video_sys_0_mm_video_bridge_s0_readdatavalid
	wire          mm_interconnect_2_video_sys_0_mm_video_bridge_s0_write;                   // mm_interconnect_2:video_sys_0_mm_video_bridge_s0_write -> video_sys_0:mm_video_bridge_s0_write
	wire   [31:0] mm_interconnect_2_video_sys_0_mm_video_bridge_s0_writedata;               // mm_interconnect_2:video_sys_0_mm_video_bridge_s0_writedata -> video_sys_0:mm_video_bridge_s0_writedata
	wire    [0:0] mm_interconnect_2_video_sys_0_mm_video_bridge_s0_burstcount;              // mm_interconnect_2:video_sys_0_mm_video_bridge_s0_burstcount -> video_sys_0:mm_video_bridge_s0_burstcount
	wire   [26:0] mm_interconnect_2_emif_bank3a_s0_axil_awaddr;                             // mm_interconnect_2:emif_bank3a_s0_axil_awaddr -> emif_bank3a:s0_axil_awaddr
	wire    [1:0] mm_interconnect_2_emif_bank3a_s0_axil_bresp;                              // emif_bank3a:s0_axil_bresp -> mm_interconnect_2:emif_bank3a_s0_axil_bresp
	wire          mm_interconnect_2_emif_bank3a_s0_axil_arready;                            // emif_bank3a:s0_axil_arready -> mm_interconnect_2:emif_bank3a_s0_axil_arready
	wire   [31:0] mm_interconnect_2_emif_bank3a_s0_axil_rdata;                              // emif_bank3a:s0_axil_rdata -> mm_interconnect_2:emif_bank3a_s0_axil_rdata
	wire    [3:0] mm_interconnect_2_emif_bank3a_s0_axil_wstrb;                              // mm_interconnect_2:emif_bank3a_s0_axil_wstrb -> emif_bank3a:s0_axil_wstrb
	wire          mm_interconnect_2_emif_bank3a_s0_axil_wready;                             // emif_bank3a:s0_axil_wready -> mm_interconnect_2:emif_bank3a_s0_axil_wready
	wire          mm_interconnect_2_emif_bank3a_s0_axil_awready;                            // emif_bank3a:s0_axil_awready -> mm_interconnect_2:emif_bank3a_s0_axil_awready
	wire          mm_interconnect_2_emif_bank3a_s0_axil_rready;                             // mm_interconnect_2:emif_bank3a_s0_axil_rready -> emif_bank3a:s0_axil_rready
	wire          mm_interconnect_2_emif_bank3a_s0_axil_bready;                             // mm_interconnect_2:emif_bank3a_s0_axil_bready -> emif_bank3a:s0_axil_bready
	wire          mm_interconnect_2_emif_bank3a_s0_axil_wvalid;                             // mm_interconnect_2:emif_bank3a_s0_axil_wvalid -> emif_bank3a:s0_axil_wvalid
	wire   [26:0] mm_interconnect_2_emif_bank3a_s0_axil_araddr;                             // mm_interconnect_2:emif_bank3a_s0_axil_araddr -> emif_bank3a:s0_axil_araddr
	wire    [2:0] mm_interconnect_2_emif_bank3a_s0_axil_arprot;                             // mm_interconnect_2:emif_bank3a_s0_axil_arprot -> emif_bank3a:s0_axil_arprot
	wire    [1:0] mm_interconnect_2_emif_bank3a_s0_axil_rresp;                              // emif_bank3a:s0_axil_rresp -> mm_interconnect_2:emif_bank3a_s0_axil_rresp
	wire    [2:0] mm_interconnect_2_emif_bank3a_s0_axil_awprot;                             // mm_interconnect_2:emif_bank3a_s0_axil_awprot -> emif_bank3a:s0_axil_awprot
	wire   [31:0] mm_interconnect_2_emif_bank3a_s0_axil_wdata;                              // mm_interconnect_2:emif_bank3a_s0_axil_wdata -> emif_bank3a:s0_axil_wdata
	wire          mm_interconnect_2_emif_bank3a_s0_axil_arvalid;                            // mm_interconnect_2:emif_bank3a_s0_axil_arvalid -> emif_bank3a:s0_axil_arvalid
	wire          mm_interconnect_2_emif_bank3a_s0_axil_bvalid;                             // emif_bank3a:s0_axil_bvalid -> mm_interconnect_2:emif_bank3a_s0_axil_bvalid
	wire          mm_interconnect_2_emif_bank3a_s0_axil_awvalid;                            // mm_interconnect_2:emif_bank3a_s0_axil_awvalid -> emif_bank3a:s0_axil_awvalid
	wire          mm_interconnect_2_emif_bank3a_s0_axil_rvalid;                             // emif_bank3a:s0_axil_rvalid -> mm_interconnect_2:emif_bank3a_s0_axil_rvalid
	wire   [31:0] bank3a_emif_master_master_readdata;                                       // mm_interconnect_3:bank3a_emif_master_master_readdata -> bank3a_emif_master:master_readdata
	wire          bank3a_emif_master_master_waitrequest;                                    // mm_interconnect_3:bank3a_emif_master_master_waitrequest -> bank3a_emif_master:master_waitrequest
	wire   [31:0] bank3a_emif_master_master_address;                                        // bank3a_emif_master:master_address -> mm_interconnect_3:bank3a_emif_master_master_address
	wire          bank3a_emif_master_master_read;                                           // bank3a_emif_master:master_read -> mm_interconnect_3:bank3a_emif_master_master_read
	wire    [3:0] bank3a_emif_master_master_byteenable;                                     // bank3a_emif_master:master_byteenable -> mm_interconnect_3:bank3a_emif_master_master_byteenable
	wire          bank3a_emif_master_master_readdatavalid;                                  // mm_interconnect_3:bank3a_emif_master_master_readdatavalid -> bank3a_emif_master:master_readdatavalid
	wire          bank3a_emif_master_master_write;                                          // bank3a_emif_master:master_write -> mm_interconnect_3:bank3a_emif_master_master_write
	wire   [31:0] bank3a_emif_master_master_writedata;                                      // bank3a_emif_master:master_writedata -> mm_interconnect_3:bank3a_emif_master_master_writedata
	wire   [63:0] mm_interconnect_3_emif_bank3a_s0_axi4_ruser;                              // emif_bank3a:s0_axi4_ruser -> mm_interconnect_3:emif_bank3a_s0_axi4_ruser
	wire   [63:0] mm_interconnect_3_emif_bank3a_s0_axi4_wuser;                              // mm_interconnect_3:emif_bank3a_s0_axi4_wuser -> emif_bank3a:s0_axi4_wuser
	wire    [1:0] mm_interconnect_3_emif_bank3a_s0_axi4_awburst;                            // mm_interconnect_3:emif_bank3a_s0_axi4_awburst -> emif_bank3a:s0_axi4_awburst
	wire   [13:0] mm_interconnect_3_emif_bank3a_s0_axi4_awuser;                             // mm_interconnect_3:emif_bank3a_s0_axi4_awuser -> emif_bank3a:s0_axi4_awuser
	wire    [7:0] mm_interconnect_3_emif_bank3a_s0_axi4_arlen;                              // mm_interconnect_3:emif_bank3a_s0_axi4_arlen -> emif_bank3a:s0_axi4_arlen
	wire    [3:0] mm_interconnect_3_emif_bank3a_s0_axi4_arqos;                              // mm_interconnect_3:emif_bank3a_s0_axi4_arqos -> emif_bank3a:s0_axi4_arqos
	wire   [31:0] mm_interconnect_3_emif_bank3a_s0_axi4_wstrb;                              // mm_interconnect_3:emif_bank3a_s0_axi4_wstrb -> emif_bank3a:s0_axi4_wstrb
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_wready;                             // emif_bank3a:s0_axi4_wready -> mm_interconnect_3:emif_bank3a_s0_axi4_wready
	wire    [6:0] mm_interconnect_3_emif_bank3a_s0_axi4_rid;                                // emif_bank3a:s0_axi4_rid -> mm_interconnect_3:emif_bank3a_s0_axi4_rid
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_rready;                             // mm_interconnect_3:emif_bank3a_s0_axi4_rready -> emif_bank3a:s0_axi4_rready
	wire    [7:0] mm_interconnect_3_emif_bank3a_s0_axi4_awlen;                              // mm_interconnect_3:emif_bank3a_s0_axi4_awlen -> emif_bank3a:s0_axi4_awlen
	wire    [3:0] mm_interconnect_3_emif_bank3a_s0_axi4_awqos;                              // mm_interconnect_3:emif_bank3a_s0_axi4_awqos -> emif_bank3a:s0_axi4_awqos
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_wvalid;                             // mm_interconnect_3:emif_bank3a_s0_axi4_wvalid -> emif_bank3a:s0_axi4_wvalid
	wire   [31:0] mm_interconnect_3_emif_bank3a_s0_axi4_araddr;                             // mm_interconnect_3:emif_bank3a_s0_axi4_araddr -> emif_bank3a:s0_axi4_araddr
	wire    [2:0] mm_interconnect_3_emif_bank3a_s0_axi4_arprot;                             // mm_interconnect_3:emif_bank3a_s0_axi4_arprot -> emif_bank3a:s0_axi4_arprot
	wire    [2:0] mm_interconnect_3_emif_bank3a_s0_axi4_awprot;                             // mm_interconnect_3:emif_bank3a_s0_axi4_awprot -> emif_bank3a:s0_axi4_awprot
	wire  [255:0] mm_interconnect_3_emif_bank3a_s0_axi4_wdata;                              // mm_interconnect_3:emif_bank3a_s0_axi4_wdata -> emif_bank3a:s0_axi4_wdata
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_arvalid;                            // mm_interconnect_3:emif_bank3a_s0_axi4_arvalid -> emif_bank3a:s0_axi4_arvalid
	wire    [6:0] mm_interconnect_3_emif_bank3a_s0_axi4_arid;                               // mm_interconnect_3:emif_bank3a_s0_axi4_arid -> emif_bank3a:s0_axi4_arid
	wire    [0:0] mm_interconnect_3_emif_bank3a_s0_axi4_arlock;                             // mm_interconnect_3:emif_bank3a_s0_axi4_arlock -> emif_bank3a:s0_axi4_arlock
	wire    [0:0] mm_interconnect_3_emif_bank3a_s0_axi4_awlock;                             // mm_interconnect_3:emif_bank3a_s0_axi4_awlock -> emif_bank3a:s0_axi4_awlock
	wire   [31:0] mm_interconnect_3_emif_bank3a_s0_axi4_awaddr;                             // mm_interconnect_3:emif_bank3a_s0_axi4_awaddr -> emif_bank3a:s0_axi4_awaddr
	wire    [1:0] mm_interconnect_3_emif_bank3a_s0_axi4_bresp;                              // emif_bank3a:s0_axi4_bresp -> mm_interconnect_3:emif_bank3a_s0_axi4_bresp
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_arready;                            // emif_bank3a:s0_axi4_arready -> mm_interconnect_3:emif_bank3a_s0_axi4_arready
	wire  [255:0] mm_interconnect_3_emif_bank3a_s0_axi4_rdata;                              // emif_bank3a:s0_axi4_rdata -> mm_interconnect_3:emif_bank3a_s0_axi4_rdata
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_awready;                            // emif_bank3a:s0_axi4_awready -> mm_interconnect_3:emif_bank3a_s0_axi4_awready
	wire    [1:0] mm_interconnect_3_emif_bank3a_s0_axi4_arburst;                            // mm_interconnect_3:emif_bank3a_s0_axi4_arburst -> emif_bank3a:s0_axi4_arburst
	wire    [2:0] mm_interconnect_3_emif_bank3a_s0_axi4_arsize;                             // mm_interconnect_3:emif_bank3a_s0_axi4_arsize -> emif_bank3a:s0_axi4_arsize
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_bready;                             // mm_interconnect_3:emif_bank3a_s0_axi4_bready -> emif_bank3a:s0_axi4_bready
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_rlast;                              // emif_bank3a:s0_axi4_rlast -> mm_interconnect_3:emif_bank3a_s0_axi4_rlast
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_wlast;                              // mm_interconnect_3:emif_bank3a_s0_axi4_wlast -> emif_bank3a:s0_axi4_wlast
	wire    [1:0] mm_interconnect_3_emif_bank3a_s0_axi4_rresp;                              // emif_bank3a:s0_axi4_rresp -> mm_interconnect_3:emif_bank3a_s0_axi4_rresp
	wire    [6:0] mm_interconnect_3_emif_bank3a_s0_axi4_awid;                               // mm_interconnect_3:emif_bank3a_s0_axi4_awid -> emif_bank3a:s0_axi4_awid
	wire    [6:0] mm_interconnect_3_emif_bank3a_s0_axi4_bid;                                // emif_bank3a:s0_axi4_bid -> mm_interconnect_3:emif_bank3a_s0_axi4_bid
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_bvalid;                             // emif_bank3a:s0_axi4_bvalid -> mm_interconnect_3:emif_bank3a_s0_axi4_bvalid
	wire    [2:0] mm_interconnect_3_emif_bank3a_s0_axi4_awsize;                             // mm_interconnect_3:emif_bank3a_s0_axi4_awsize -> emif_bank3a:s0_axi4_awsize
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_awvalid;                            // mm_interconnect_3:emif_bank3a_s0_axi4_awvalid -> emif_bank3a:s0_axi4_awvalid
	wire   [13:0] mm_interconnect_3_emif_bank3a_s0_axi4_aruser;                             // mm_interconnect_3:emif_bank3a_s0_axi4_aruser -> emif_bank3a:s0_axi4_aruser
	wire          mm_interconnect_3_emif_bank3a_s0_axi4_rvalid;                             // emif_bank3a:s0_axi4_rvalid -> mm_interconnect_3:emif_bank3a_s0_axi4_rvalid
	wire          irq_mapper_receiver0_irq;                                                 // peripheral_sys_0:dipsw_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                 // video_sys_0:hdmi_dmac_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                 // peripheral_sys_0:jtag_uart_irq_irq -> irq_mapper:receiver2_irq
	wire          irq_mapper_receiver3_irq;                                                 // peripheral_sys_0:pb_irq_irq -> irq_mapper:receiver3_irq
	wire   [62:0] agilex_5_soc_fpga2hps_interrupt_irq;                                      // irq_mapper:sender_irq -> agilex_5_soc:fpga2hps_interrupt_irq
	wire          rst_controller_reset_out_reset;                                           // rst_controller:reset_out -> emif_bank3a:core_init_n_0
	wire          agilex_5_soc_h2f_cold_reset_reset;                                        // agilex_5_soc:h2f_cold_reset_reset_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_007:reset_in0]
	wire          agilex_5_soc_h2f_reset_reset;                                             // agilex_5_soc:h2f_reset_reset_n -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_007:reset_in1]
	wire          rst_controller_001_reset_out_reset;                                       // rst_controller_001:reset_out -> emif_bank3a:s0_axil_rst_n
	wire          rst_controller_002_reset_out_reset;                                       // rst_controller_002:reset_out -> fpga_only_master:clk_reset_reset
	wire          fpga_only_master_master_reset_reset;                                      // fpga_only_master:master_reset_reset -> [rst_controller_002:reset_in0, rst_controller_006:reset_in0]
	wire          rst_controller_003_reset_out_reset;                                       // rst_controller_003:reset_out -> onchip_sram:reset
	wire          rst_controller_004_reset_out_reset;                                       // rst_controller_004:reset_out -> [mm_interconnect_0:f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_1:agilex_5_soc_hps2fpga_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:peripheral_sys_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:agilex_5_soc_lwhps2fpga_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_2:video_sys_0_reset_reset_bridge_in_reset_reset, mm_interconnect_3:bank3a_emif_master_master_translator_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_005_reset_out_reset;                                       // rst_controller_005:reset_out -> [mm_interconnect_1:onchip_sram_axi_s1_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:onchip_sram_reset1_reset_bridge_in_reset_reset]
	wire          rst_controller_006_reset_out_reset;                                       // rst_controller_006:reset_out -> [mm_interconnect_1:crosser_002_in_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:fpga_only_master_master_translator_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_007_reset_out_reset;                                       // rst_controller_007:reset_out -> mm_interconnect_2:emif_bank3a_s0_axil_agent_reset_sink_reset_bridge_in_reset_reset
	wire          rst_controller_008_reset_out_reset;                                       // rst_controller_008:reset_out -> mm_interconnect_3:emif_bank3a_s0_axi4_translator_clk_reset_reset_bridge_in_reset_reset
	wire          emif_bank3a_usr_rst_n_0_reset;                                            // emif_bank3a:usr_rst_n_0 -> rst_controller_008:reset_in0

	ghrd_hps_system_intel_agilex_5_soc_0 agilex_5_soc (
		.h2f_reset_reset_n                  (agilex_5_soc_h2f_reset_reset),                    //  output,    width = 1,                h2f_reset.reset_n
		.hps2fpga_axi_clock_clk             (agilex_5_soc_h2f_user1_clk_clk),                  //   input,    width = 1,       hps2fpga_axi_clock.clk
		.hps2fpga_axi_reset_reset_n         (~reset_in_out_reset_reset),                       //   input,    width = 1,       hps2fpga_axi_reset.reset_n
		.hps2fpga_awid                      (agilex_5_soc_hps2fpga_awid),                      //  output,    width = 4,                 hps2fpga.awid
		.hps2fpga_awaddr                    (agilex_5_soc_hps2fpga_awaddr),                    //  output,   width = 32,                         .awaddr
		.hps2fpga_awlen                     (agilex_5_soc_hps2fpga_awlen),                     //  output,    width = 8,                         .awlen
		.hps2fpga_awsize                    (agilex_5_soc_hps2fpga_awsize),                    //  output,    width = 3,                         .awsize
		.hps2fpga_awburst                   (agilex_5_soc_hps2fpga_awburst),                   //  output,    width = 2,                         .awburst
		.hps2fpga_awlock                    (agilex_5_soc_hps2fpga_awlock),                    //  output,    width = 1,                         .awlock
		.hps2fpga_awcache                   (agilex_5_soc_hps2fpga_awcache),                   //  output,    width = 4,                         .awcache
		.hps2fpga_awprot                    (agilex_5_soc_hps2fpga_awprot),                    //  output,    width = 3,                         .awprot
		.hps2fpga_awvalid                   (agilex_5_soc_hps2fpga_awvalid),                   //  output,    width = 1,                         .awvalid
		.hps2fpga_awready                   (agilex_5_soc_hps2fpga_awready),                   //   input,    width = 1,                         .awready
		.hps2fpga_wdata                     (agilex_5_soc_hps2fpga_wdata),                     //  output,   width = 32,                         .wdata
		.hps2fpga_wstrb                     (agilex_5_soc_hps2fpga_wstrb),                     //  output,    width = 4,                         .wstrb
		.hps2fpga_wlast                     (agilex_5_soc_hps2fpga_wlast),                     //  output,    width = 1,                         .wlast
		.hps2fpga_wvalid                    (agilex_5_soc_hps2fpga_wvalid),                    //  output,    width = 1,                         .wvalid
		.hps2fpga_wready                    (agilex_5_soc_hps2fpga_wready),                    //   input,    width = 1,                         .wready
		.hps2fpga_bid                       (agilex_5_soc_hps2fpga_bid),                       //   input,    width = 4,                         .bid
		.hps2fpga_bresp                     (agilex_5_soc_hps2fpga_bresp),                     //   input,    width = 2,                         .bresp
		.hps2fpga_bvalid                    (agilex_5_soc_hps2fpga_bvalid),                    //   input,    width = 1,                         .bvalid
		.hps2fpga_bready                    (agilex_5_soc_hps2fpga_bready),                    //  output,    width = 1,                         .bready
		.hps2fpga_arid                      (agilex_5_soc_hps2fpga_arid),                      //  output,    width = 4,                         .arid
		.hps2fpga_araddr                    (agilex_5_soc_hps2fpga_araddr),                    //  output,   width = 32,                         .araddr
		.hps2fpga_arlen                     (agilex_5_soc_hps2fpga_arlen),                     //  output,    width = 8,                         .arlen
		.hps2fpga_arsize                    (agilex_5_soc_hps2fpga_arsize),                    //  output,    width = 3,                         .arsize
		.hps2fpga_arburst                   (agilex_5_soc_hps2fpga_arburst),                   //  output,    width = 2,                         .arburst
		.hps2fpga_arlock                    (agilex_5_soc_hps2fpga_arlock),                    //  output,    width = 1,                         .arlock
		.hps2fpga_arcache                   (agilex_5_soc_hps2fpga_arcache),                   //  output,    width = 4,                         .arcache
		.hps2fpga_arprot                    (agilex_5_soc_hps2fpga_arprot),                    //  output,    width = 3,                         .arprot
		.hps2fpga_arvalid                   (agilex_5_soc_hps2fpga_arvalid),                   //  output,    width = 1,                         .arvalid
		.hps2fpga_arready                   (agilex_5_soc_hps2fpga_arready),                   //   input,    width = 1,                         .arready
		.hps2fpga_rid                       (agilex_5_soc_hps2fpga_rid),                       //   input,    width = 4,                         .rid
		.hps2fpga_rdata                     (agilex_5_soc_hps2fpga_rdata),                     //   input,   width = 32,                         .rdata
		.hps2fpga_rresp                     (agilex_5_soc_hps2fpga_rresp),                     //   input,    width = 2,                         .rresp
		.hps2fpga_rlast                     (agilex_5_soc_hps2fpga_rlast),                     //   input,    width = 1,                         .rlast
		.hps2fpga_rvalid                    (agilex_5_soc_hps2fpga_rvalid),                    //   input,    width = 1,                         .rvalid
		.hps2fpga_rready                    (agilex_5_soc_hps2fpga_rready),                    //  output,    width = 1,                         .rready
		.lwhps2fpga_axi_clock_clk           (agilex_5_soc_h2f_user1_clk_clk),                  //   input,    width = 1,     lwhps2fpga_axi_clock.clk
		.lwhps2fpga_axi_reset_reset_n       (~reset_in_out_reset_reset),                       //   input,    width = 1,     lwhps2fpga_axi_reset.reset_n
		.lwhps2fpga_awid                    (agilex_5_soc_lwhps2fpga_awid),                    //  output,    width = 4,               lwhps2fpga.awid
		.lwhps2fpga_awaddr                  (agilex_5_soc_lwhps2fpga_awaddr),                  //  output,   width = 29,                         .awaddr
		.lwhps2fpga_awlen                   (agilex_5_soc_lwhps2fpga_awlen),                   //  output,    width = 8,                         .awlen
		.lwhps2fpga_awsize                  (agilex_5_soc_lwhps2fpga_awsize),                  //  output,    width = 3,                         .awsize
		.lwhps2fpga_awburst                 (agilex_5_soc_lwhps2fpga_awburst),                 //  output,    width = 2,                         .awburst
		.lwhps2fpga_awlock                  (agilex_5_soc_lwhps2fpga_awlock),                  //  output,    width = 1,                         .awlock
		.lwhps2fpga_awcache                 (agilex_5_soc_lwhps2fpga_awcache),                 //  output,    width = 4,                         .awcache
		.lwhps2fpga_awprot                  (agilex_5_soc_lwhps2fpga_awprot),                  //  output,    width = 3,                         .awprot
		.lwhps2fpga_awvalid                 (agilex_5_soc_lwhps2fpga_awvalid),                 //  output,    width = 1,                         .awvalid
		.lwhps2fpga_awready                 (agilex_5_soc_lwhps2fpga_awready),                 //   input,    width = 1,                         .awready
		.lwhps2fpga_wdata                   (agilex_5_soc_lwhps2fpga_wdata),                   //  output,   width = 32,                         .wdata
		.lwhps2fpga_wstrb                   (agilex_5_soc_lwhps2fpga_wstrb),                   //  output,    width = 4,                         .wstrb
		.lwhps2fpga_wlast                   (agilex_5_soc_lwhps2fpga_wlast),                   //  output,    width = 1,                         .wlast
		.lwhps2fpga_wvalid                  (agilex_5_soc_lwhps2fpga_wvalid),                  //  output,    width = 1,                         .wvalid
		.lwhps2fpga_wready                  (agilex_5_soc_lwhps2fpga_wready),                  //   input,    width = 1,                         .wready
		.lwhps2fpga_bid                     (agilex_5_soc_lwhps2fpga_bid),                     //   input,    width = 4,                         .bid
		.lwhps2fpga_bresp                   (agilex_5_soc_lwhps2fpga_bresp),                   //   input,    width = 2,                         .bresp
		.lwhps2fpga_bvalid                  (agilex_5_soc_lwhps2fpga_bvalid),                  //   input,    width = 1,                         .bvalid
		.lwhps2fpga_bready                  (agilex_5_soc_lwhps2fpga_bready),                  //  output,    width = 1,                         .bready
		.lwhps2fpga_arid                    (agilex_5_soc_lwhps2fpga_arid),                    //  output,    width = 4,                         .arid
		.lwhps2fpga_araddr                  (agilex_5_soc_lwhps2fpga_araddr),                  //  output,   width = 29,                         .araddr
		.lwhps2fpga_arlen                   (agilex_5_soc_lwhps2fpga_arlen),                   //  output,    width = 8,                         .arlen
		.lwhps2fpga_arsize                  (agilex_5_soc_lwhps2fpga_arsize),                  //  output,    width = 3,                         .arsize
		.lwhps2fpga_arburst                 (agilex_5_soc_lwhps2fpga_arburst),                 //  output,    width = 2,                         .arburst
		.lwhps2fpga_arlock                  (agilex_5_soc_lwhps2fpga_arlock),                  //  output,    width = 1,                         .arlock
		.lwhps2fpga_arcache                 (agilex_5_soc_lwhps2fpga_arcache),                 //  output,    width = 4,                         .arcache
		.lwhps2fpga_arprot                  (agilex_5_soc_lwhps2fpga_arprot),                  //  output,    width = 3,                         .arprot
		.lwhps2fpga_arvalid                 (agilex_5_soc_lwhps2fpga_arvalid),                 //  output,    width = 1,                         .arvalid
		.lwhps2fpga_arready                 (agilex_5_soc_lwhps2fpga_arready),                 //   input,    width = 1,                         .arready
		.lwhps2fpga_rid                     (agilex_5_soc_lwhps2fpga_rid),                     //   input,    width = 4,                         .rid
		.lwhps2fpga_rdata                   (agilex_5_soc_lwhps2fpga_rdata),                   //   input,   width = 32,                         .rdata
		.lwhps2fpga_rresp                   (agilex_5_soc_lwhps2fpga_rresp),                   //   input,    width = 2,                         .rresp
		.lwhps2fpga_rlast                   (agilex_5_soc_lwhps2fpga_rlast),                   //   input,    width = 1,                         .rlast
		.lwhps2fpga_rvalid                  (agilex_5_soc_lwhps2fpga_rvalid),                  //   input,    width = 1,                         .rvalid
		.lwhps2fpga_rready                  (agilex_5_soc_lwhps2fpga_rready),                  //  output,    width = 1,                         .rready
		.emac_ptp_clk_clk                   (agilex_5_soc_h2f_user0_clk_clk),                  //   input,    width = 1,             emac_ptp_clk.clk
		.emac_timestamp_clk_clk             (agilex_5_soc_h2f_user0_clk_clk),                  //   input,    width = 1,       emac_timestamp_clk.clk
		.emac_timestamp_data_data_in        (),                                                //   input,   width = 64,      emac_timestamp_data.data_in
		.emac0_mdio_mac_mdc                 (emac0_mdio_mac_mdc),                              //  output,    width = 1,               emac0_mdio.mac_mdc
		.emac0_mdio_mac_mdi                 (emac0_mdio_mac_mdi),                              //   input,    width = 1,                         .mac_mdi
		.emac0_mdio_mac_mdo                 (emac0_mdio_mac_mdo),                              //  output,    width = 1,                         .mac_mdo
		.emac0_mdio_mac_mdoe                (emac0_mdio_mac_mdoe),                             //  output,    width = 1,                         .mac_mdoe
		.emac0_app_rst_reset_n              (emac0_app_rst_reset_n),                           //  output,    width = 1,            emac0_app_rst.reset_n
		.emac0_mac_tx_clk_o                 (emac0_mac_tx_clk_o),                              //  output,    width = 1,                    emac0.mac_tx_clk_o
		.emac0_mac_tx_clk_i                 (emac0_mac_tx_clk_i),                              //   input,    width = 1,                         .mac_tx_clk_i
		.emac0_mac_rx_clk                   (emac0_mac_rx_clk),                                //   input,    width = 1,                         .mac_rx_clk
		.emac0_mac_rst_tx_n                 (emac0_mac_rst_tx_n),                              //  output,    width = 1,                         .mac_rst_tx_n
		.emac0_mac_rst_rx_n                 (emac0_mac_rst_rx_n),                              //  output,    width = 1,                         .mac_rst_rx_n
		.emac0_mac_txen                     (emac0_mac_txen),                                  //  output,    width = 1,                         .mac_txen
		.emac0_mac_txer                     (emac0_mac_txer),                                  //  output,    width = 1,                         .mac_txer
		.emac0_mac_rxdv                     (emac0_mac_rxdv),                                  //   input,    width = 1,                         .mac_rxdv
		.emac0_mac_rxer                     (emac0_mac_rxer),                                  //   input,    width = 1,                         .mac_rxer
		.emac0_mac_rxd                      (emac0_mac_rxd),                                   //   input,    width = 8,                         .mac_rxd
		.emac0_mac_col                      (emac0_mac_col),                                   //   input,    width = 1,                         .mac_col
		.emac0_mac_crs                      (emac0_mac_crs),                                   //   input,    width = 1,                         .mac_crs
		.emac0_mac_speed                    (emac0_mac_speed),                                 //  output,    width = 3,                         .mac_speed
		.emac0_mac_txd_o                    (emac0_mac_txd_o),                                 //  output,    width = 8,                         .mac_txd_o
		.emac2_app_rst_reset_n              (emac2_app_rst_reset_n),                           //  output,    width = 1,            emac2_app_rst.reset_n
		.spim0_miso_i                       (spim0_miso_i),                                    //   input,    width = 1,                    spim0.miso_i
		.spim0_mosi_o                       (spim0_mosi_o),                                    //  output,    width = 1,                         .mosi_o
		.spim0_mosi_oe                      (spim0_mosi_oe),                                   //  output,    width = 1,                         .mosi_oe
		.spim0_ss_in_n                      (spim0_ss_in_n),                                   //   input,    width = 1,                         .ss_in_n
		.spim0_ss0_n_o                      (spim0_ss0_n_o),                                   //  output,    width = 1,                         .ss0_n_o
		.spim0_ss1_n_o                      (spim0_ss1_n_o),                                   //  output,    width = 1,                         .ss1_n_o
		.spim0_ss2_n_o                      (spim0_ss2_n_o),                                   //  output,    width = 1,                         .ss2_n_o
		.spim0_ss3_n_o                      (spim0_ss3_n_o),                                   //  output,    width = 1,                         .ss3_n_o
		.spim0_sclk_out_clk                 (spim0_sclk_out_clk),                              //  output,    width = 1,           spim0_sclk_out.clk
		.I2C1_scl_i_clk                     (i2c1_scl_i_clk),                                  //   input,    width = 1,               I2C1_scl_i.clk
		.I2C1_scl_oe_clk                    (i2c1_scl_oe_clk),                                 //  output,    width = 1,              I2C1_scl_oe.clk
		.I2C1_sda_i                         (i2c1_sda_i),                                      //   input,    width = 1,                     I2C1.sda_i
		.I2C1_sda_oe                        (i2c1_sda_oe),                                     //  output,    width = 1,                         .sda_oe
		.h2f_user0_clk_clk                  (agilex_5_soc_h2f_user0_clk_clk),                  //  output,    width = 1,            h2f_user0_clk.clk
		.h2f_user1_clk_clk                  (agilex_5_soc_h2f_user1_clk_clk),                  //  output,    width = 1,            h2f_user1_clk.clk
		.h2f_warm_reset_handshake_reset_req (),                                                //  output,    width = 1, h2f_warm_reset_handshake.reset_req
		.h2f_warm_reset_handshake_reset_ack (),                                                //   input,    width = 1,                         .reset_ack
		.h2f_cold_reset_reset_n             (agilex_5_soc_h2f_cold_reset_reset),               //  output,    width = 1,           h2f_cold_reset.reset_n
		.hps_io_hps_osc_clk                 (hps_io_hps_osc_clk),                              //   input,    width = 1,                   hps_io.hps_osc_clk
		.hps_io_sdmmc_data0                 (hps_io_sdmmc_data0),                              //   inout,    width = 1,                         .sdmmc_data0
		.hps_io_sdmmc_data1                 (hps_io_sdmmc_data1),                              //   inout,    width = 1,                         .sdmmc_data1
		.hps_io_sdmmc_cclk                  (hps_io_sdmmc_cclk),                               //  output,    width = 1,                         .sdmmc_cclk
		.hps_io_sdmmc_data2                 (hps_io_sdmmc_data2),                              //   inout,    width = 1,                         .sdmmc_data2
		.hps_io_sdmmc_data3                 (hps_io_sdmmc_data3),                              //   inout,    width = 1,                         .sdmmc_data3
		.hps_io_sdmmc_cmd                   (hps_io_sdmmc_cmd),                                //   inout,    width = 1,                         .sdmmc_cmd
		.hps_io_usb1_clk                    (hps_io_usb1_clk),                                 //   input,    width = 1,                         .usb1_clk
		.hps_io_usb1_stp                    (hps_io_usb1_stp),                                 //  output,    width = 1,                         .usb1_stp
		.hps_io_usb1_dir                    (hps_io_usb1_dir),                                 //   input,    width = 1,                         .usb1_dir
		.hps_io_usb1_data0                  (hps_io_usb1_data0),                               //   inout,    width = 1,                         .usb1_data0
		.hps_io_usb1_data1                  (hps_io_usb1_data1),                               //   inout,    width = 1,                         .usb1_data1
		.hps_io_usb1_nxr                    (hps_io_usb1_nxr),                                 //   input,    width = 1,                         .usb1_nxr
		.hps_io_usb1_data2                  (hps_io_usb1_data2),                               //   inout,    width = 1,                         .usb1_data2
		.hps_io_usb1_data3                  (hps_io_usb1_data3),                               //   inout,    width = 1,                         .usb1_data3
		.hps_io_usb1_data4                  (hps_io_usb1_data4),                               //   inout,    width = 1,                         .usb1_data4
		.hps_io_usb1_data5                  (hps_io_usb1_data5),                               //   inout,    width = 1,                         .usb1_data5
		.hps_io_usb1_data6                  (hps_io_usb1_data6),                               //   inout,    width = 1,                         .usb1_data6
		.hps_io_usb1_data7                  (hps_io_usb1_data7),                               //   inout,    width = 1,                         .usb1_data7
		.hps_io_emac2_tx_clk                (hps_io_emac2_tx_clk),                             //  output,    width = 1,                         .emac2_tx_clk
		.hps_io_emac2_tx_ctl                (hps_io_emac2_tx_ctl),                             //  output,    width = 1,                         .emac2_tx_ctl
		.hps_io_emac2_rx_clk                (hps_io_emac2_rx_clk),                             //   input,    width = 1,                         .emac2_rx_clk
		.hps_io_emac2_rx_ctl                (hps_io_emac2_rx_ctl),                             //   input,    width = 1,                         .emac2_rx_ctl
		.hps_io_emac2_txd0                  (hps_io_emac2_txd0),                               //  output,    width = 1,                         .emac2_txd0
		.hps_io_emac2_txd1                  (hps_io_emac2_txd1),                               //  output,    width = 1,                         .emac2_txd1
		.hps_io_emac2_rxd0                  (hps_io_emac2_rxd0),                               //   input,    width = 1,                         .emac2_rxd0
		.hps_io_emac2_rxd1                  (hps_io_emac2_rxd1),                               //   input,    width = 1,                         .emac2_rxd1
		.hps_io_emac2_txd2                  (hps_io_emac2_txd2),                               //  output,    width = 1,                         .emac2_txd2
		.hps_io_emac2_txd3                  (hps_io_emac2_txd3),                               //  output,    width = 1,                         .emac2_txd3
		.hps_io_emac2_rxd2                  (hps_io_emac2_rxd2),                               //   input,    width = 1,                         .emac2_rxd2
		.hps_io_emac2_rxd3                  (hps_io_emac2_rxd3),                               //   input,    width = 1,                         .emac2_rxd3
		.hps_io_mdio2_mdio                  (hps_io_mdio2_mdio),                               //   inout,    width = 1,                         .mdio2_mdio
		.hps_io_mdio2_mdc                   (hps_io_mdio2_mdc),                                //  output,    width = 1,                         .mdio2_mdc
		.hps_io_uart0_tx                    (hps_io_uart0_tx),                                 //  output,    width = 1,                         .uart0_tx
		.hps_io_uart0_rx                    (hps_io_uart0_rx),                                 //   input,    width = 1,                         .uart0_rx
		.hps_io_i2c0_sda                    (hps_io_i2c0_sda),                                 //   inout,    width = 1,                         .i2c0_sda
		.hps_io_i2c0_scl                    (hps_io_i2c0_scl),                                 //   inout,    width = 1,                         .i2c0_scl
		.hps_io_gpio6                       (hps_io_gpio6),                                    //   inout,    width = 1,                         .gpio6
		.hps_io_gpio7                       (hps_io_gpio7),                                    //   inout,    width = 1,                         .gpio7
		.hps_io_gpio8                       (hps_io_gpio8),                                    //   inout,    width = 1,                         .gpio8
		.hps_io_gpio9                       (hps_io_gpio9),                                    //   inout,    width = 1,                         .gpio9
		.hps_io_gpio10                      (hps_io_gpio10),                                   //   inout,    width = 1,                         .gpio10
		.hps_io_gpio11                      (hps_io_gpio11),                                   //   inout,    width = 1,                         .gpio11
		.hps_io_gpio28                      (hps_io_gpio28),                                   //   inout,    width = 1,                         .gpio28
		.hps_io_gpio34                      (hps_io_gpio34),                                   //   inout,    width = 1,                         .gpio34
		.hps_io_gpio35                      (hps_io_gpio35),                                   //   inout,    width = 1,                         .gpio35
		.usb31_io_vbus_det                  (usb31_io_vbus_det),                               //   input,    width = 1,                 usb31_io.vbus_det
		.usb31_io_flt_bar                   (usb31_io_flt_bar),                                //   input,    width = 1,                         .flt_bar
		.usb31_io_usb_ctrl                  (usb31_io_usb_ctrl),                               //  output,    width = 2,                         .usb_ctrl
		.usb31_io_usb31_id                  (usb31_io_usb31_id),                               //   input,    width = 1,                         .usb31_id
		.fpga2hps_interrupt_irq             (agilex_5_soc_fpga2hps_interrupt_irq),             //   input,   width = 63,       fpga2hps_interrupt.irq
		.f2sdram_axi_clock_clk              (agilex_5_soc_h2f_user1_clk_clk),                  //   input,    width = 1,        f2sdram_axi_clock.clk
		.f2sdram_axi_reset_reset_n          (~reset_in_out_reset_reset),                       //   input,    width = 1,        f2sdram_axi_reset.reset_n
		.f2sdram_araddr                     (mm_interconnect_0_agilex_5_soc_f2sdram_araddr),   //   input,   width = 32,                  f2sdram.araddr
		.f2sdram_arburst                    (mm_interconnect_0_agilex_5_soc_f2sdram_arburst),  //   input,    width = 2,                         .arburst
		.f2sdram_arcache                    (mm_interconnect_0_agilex_5_soc_f2sdram_arcache),  //   input,    width = 4,                         .arcache
		.f2sdram_arid                       (mm_interconnect_0_agilex_5_soc_f2sdram_arid),     //   input,    width = 5,                         .arid
		.f2sdram_arlen                      (mm_interconnect_0_agilex_5_soc_f2sdram_arlen),    //   input,    width = 8,                         .arlen
		.f2sdram_arlock                     (mm_interconnect_0_agilex_5_soc_f2sdram_arlock),   //   input,    width = 1,                         .arlock
		.f2sdram_arprot                     (mm_interconnect_0_agilex_5_soc_f2sdram_arprot),   //   input,    width = 3,                         .arprot
		.f2sdram_arqos                      (mm_interconnect_0_agilex_5_soc_f2sdram_arqos),    //   input,    width = 4,                         .arqos
		.f2sdram_arready                    (mm_interconnect_0_agilex_5_soc_f2sdram_arready),  //  output,    width = 1,                         .arready
		.f2sdram_arsize                     (mm_interconnect_0_agilex_5_soc_f2sdram_arsize),   //   input,    width = 3,                         .arsize
		.f2sdram_arvalid                    (mm_interconnect_0_agilex_5_soc_f2sdram_arvalid),  //   input,    width = 1,                         .arvalid
		.f2sdram_awaddr                     (mm_interconnect_0_agilex_5_soc_f2sdram_awaddr),   //   input,   width = 32,                         .awaddr
		.f2sdram_awburst                    (mm_interconnect_0_agilex_5_soc_f2sdram_awburst),  //   input,    width = 2,                         .awburst
		.f2sdram_awcache                    (mm_interconnect_0_agilex_5_soc_f2sdram_awcache),  //   input,    width = 4,                         .awcache
		.f2sdram_awid                       (mm_interconnect_0_agilex_5_soc_f2sdram_awid),     //   input,    width = 5,                         .awid
		.f2sdram_awlen                      (mm_interconnect_0_agilex_5_soc_f2sdram_awlen),    //   input,    width = 8,                         .awlen
		.f2sdram_awlock                     (mm_interconnect_0_agilex_5_soc_f2sdram_awlock),   //   input,    width = 1,                         .awlock
		.f2sdram_awprot                     (mm_interconnect_0_agilex_5_soc_f2sdram_awprot),   //   input,    width = 3,                         .awprot
		.f2sdram_awqos                      (mm_interconnect_0_agilex_5_soc_f2sdram_awqos),    //   input,    width = 4,                         .awqos
		.f2sdram_awready                    (mm_interconnect_0_agilex_5_soc_f2sdram_awready),  //  output,    width = 1,                         .awready
		.f2sdram_awsize                     (mm_interconnect_0_agilex_5_soc_f2sdram_awsize),   //   input,    width = 3,                         .awsize
		.f2sdram_awvalid                    (mm_interconnect_0_agilex_5_soc_f2sdram_awvalid),  //   input,    width = 1,                         .awvalid
		.f2sdram_bid                        (mm_interconnect_0_agilex_5_soc_f2sdram_bid),      //  output,    width = 5,                         .bid
		.f2sdram_bready                     (mm_interconnect_0_agilex_5_soc_f2sdram_bready),   //   input,    width = 1,                         .bready
		.f2sdram_bresp                      (mm_interconnect_0_agilex_5_soc_f2sdram_bresp),    //  output,    width = 2,                         .bresp
		.f2sdram_bvalid                     (mm_interconnect_0_agilex_5_soc_f2sdram_bvalid),   //  output,    width = 1,                         .bvalid
		.f2sdram_rdata                      (mm_interconnect_0_agilex_5_soc_f2sdram_rdata),    //  output,   width = 64,                         .rdata
		.f2sdram_rid                        (mm_interconnect_0_agilex_5_soc_f2sdram_rid),      //  output,    width = 5,                         .rid
		.f2sdram_rlast                      (mm_interconnect_0_agilex_5_soc_f2sdram_rlast),    //  output,    width = 1,                         .rlast
		.f2sdram_rready                     (mm_interconnect_0_agilex_5_soc_f2sdram_rready),   //   input,    width = 1,                         .rready
		.f2sdram_rresp                      (mm_interconnect_0_agilex_5_soc_f2sdram_rresp),    //  output,    width = 2,                         .rresp
		.f2sdram_rvalid                     (mm_interconnect_0_agilex_5_soc_f2sdram_rvalid),   //  output,    width = 1,                         .rvalid
		.f2sdram_wdata                      (mm_interconnect_0_agilex_5_soc_f2sdram_wdata),    //   input,   width = 64,                         .wdata
		.f2sdram_wlast                      (mm_interconnect_0_agilex_5_soc_f2sdram_wlast),    //   input,    width = 1,                         .wlast
		.f2sdram_wready                     (mm_interconnect_0_agilex_5_soc_f2sdram_wready),   //  output,    width = 1,                         .wready
		.f2sdram_wstrb                      (mm_interconnect_0_agilex_5_soc_f2sdram_wstrb),    //   input,    width = 8,                         .wstrb
		.f2sdram_wvalid                     (mm_interconnect_0_agilex_5_soc_f2sdram_wvalid),   //   input,    width = 1,                         .wvalid
		.f2sdram_aruser                     (mm_interconnect_0_agilex_5_soc_f2sdram_aruser),   //   input,    width = 8,                         .aruser
		.f2sdram_awuser                     (mm_interconnect_0_agilex_5_soc_f2sdram_awuser),   //   input,    width = 8,                         .awuser
		.f2sdram_wuser                      (mm_interconnect_0_agilex_5_soc_f2sdram_wuser),    //   input,    width = 8,                         .wuser
		.f2sdram_buser                      (mm_interconnect_0_agilex_5_soc_f2sdram_buser),    //  output,    width = 8,                         .buser
		.f2sdram_arregion                   (mm_interconnect_0_agilex_5_soc_f2sdram_arregion), //   input,    width = 4,                         .arregion
		.f2sdram_ruser                      (mm_interconnect_0_agilex_5_soc_f2sdram_ruser),    //  output,    width = 8,                         .ruser
		.f2sdram_awregion                   (mm_interconnect_0_agilex_5_soc_f2sdram_awregion), //   input,    width = 4,                         .awregion
		.fpga2hps_clock_clk                 (agilex_5_soc_h2f_user1_clk_clk),                  //   input,    width = 1,           fpga2hps_clock.clk
		.fpga2hps_reset_reset_n             (~reset_in_out_reset_reset),                       //   input,    width = 1,           fpga2hps_reset.reset_n
		.fpga2hps_awid                      (),                                                //   input,    width = 5,                 fpga2hps.awid
		.fpga2hps_awaddr                    (),                                                //   input,   width = 31,                         .awaddr
		.fpga2hps_awlen                     (),                                                //   input,    width = 8,                         .awlen
		.fpga2hps_awsize                    (),                                                //   input,    width = 3,                         .awsize
		.fpga2hps_arsize                    (),                                                //   input,    width = 3,                         .arsize
		.fpga2hps_awburst                   (),                                                //   input,    width = 2,                         .awburst
		.fpga2hps_awlock                    (),                                                //   input,    width = 1,                         .awlock
		.fpga2hps_awcache                   (),                                                //   input,    width = 4,                         .awcache
		.fpga2hps_awprot                    (),                                                //   input,    width = 3,                         .awprot
		.fpga2hps_awqos                     (),                                                //   input,    width = 4,                         .awqos
		.fpga2hps_awvalid                   (),                                                //   input,    width = 1,                         .awvalid
		.fpga2hps_awready                   (),                                                //  output,    width = 1,                         .awready
		.fpga2hps_wdata                     (),                                                //   input,  width = 256,                         .wdata
		.fpga2hps_wstrb                     (),                                                //   input,   width = 32,                         .wstrb
		.fpga2hps_wlast                     (),                                                //   input,    width = 1,                         .wlast
		.fpga2hps_wvalid                    (),                                                //   input,    width = 1,                         .wvalid
		.fpga2hps_wready                    (),                                                //  output,    width = 1,                         .wready
		.fpga2hps_bid                       (),                                                //  output,    width = 5,                         .bid
		.fpga2hps_bresp                     (),                                                //  output,    width = 2,                         .bresp
		.fpga2hps_bvalid                    (),                                                //  output,    width = 1,                         .bvalid
		.fpga2hps_bready                    (),                                                //   input,    width = 1,                         .bready
		.fpga2hps_arid                      (),                                                //   input,    width = 5,                         .arid
		.fpga2hps_araddr                    (),                                                //   input,   width = 31,                         .araddr
		.fpga2hps_arlen                     (),                                                //   input,    width = 8,                         .arlen
		.fpga2hps_arburst                   (),                                                //   input,    width = 2,                         .arburst
		.fpga2hps_arlock                    (),                                                //   input,    width = 1,                         .arlock
		.fpga2hps_arcache                   (),                                                //   input,    width = 4,                         .arcache
		.fpga2hps_arprot                    (),                                                //   input,    width = 3,                         .arprot
		.fpga2hps_arqos                     (),                                                //   input,    width = 4,                         .arqos
		.fpga2hps_arvalid                   (),                                                //   input,    width = 1,                         .arvalid
		.fpga2hps_arready                   (),                                                //  output,    width = 1,                         .arready
		.fpga2hps_rid                       (),                                                //  output,    width = 5,                         .rid
		.fpga2hps_rdata                     (),                                                //  output,  width = 256,                         .rdata
		.fpga2hps_rresp                     (),                                                //  output,    width = 2,                         .rresp
		.fpga2hps_rlast                     (),                                                //  output,    width = 1,                         .rlast
		.fpga2hps_rvalid                    (),                                                //  output,    width = 1,                         .rvalid
		.fpga2hps_rready                    (),                                                //   input,    width = 1,                         .rready
		.fpga2hps_aruser                    (),                                                //   input,    width = 8,                         .aruser
		.fpga2hps_awuser                    (),                                                //   input,    width = 8,                         .awuser
		.fpga2hps_arregion                  (),                                                //   input,    width = 4,                         .arregion
		.fpga2hps_awregion                  (),                                                //   input,    width = 4,                         .awregion
		.fpga2hps_wuser                     (),                                                //   input,    width = 8,                         .wuser
		.fpga2hps_buser                     (),                                                //  output,    width = 8,                         .buser
		.fpga2hps_ruser                     ()                                                 //  output,    width = 8,                         .ruser
	);

	ghrd_hps_system_master_0 bank3a_emif_master (
		.clk_clk              (agilex_5_soc_h2f_user1_clk_clk),          //   input,   width = 1,          clk.clk
		.clk_reset_reset      (reset_in_out_reset_reset),                //   input,   width = 1,    clk_reset.reset
		.master_reset_reset   (),                                        //  output,   width = 1, master_reset.reset
		.master_address       (bank3a_emif_master_master_address),       //  output,  width = 32,       master.address
		.master_readdata      (bank3a_emif_master_master_readdata),      //   input,  width = 32,             .readdata
		.master_read          (bank3a_emif_master_master_read),          //  output,   width = 1,             .read
		.master_write         (bank3a_emif_master_master_write),         //  output,   width = 1,             .write
		.master_writedata     (bank3a_emif_master_master_writedata),     //  output,  width = 32,             .writedata
		.master_waitrequest   (bank3a_emif_master_master_waitrequest),   //   input,   width = 1,             .waitrequest
		.master_readdatavalid (bank3a_emif_master_master_readdatavalid), //   input,   width = 1,             .readdatavalid
		.master_byteenable    (bank3a_emif_master_master_byteenable)     //  output,   width = 4,             .byteenable
	);

	emif_ph2_1 emif_bank3a (
		.ref_clk_0       (bank3a_lpddr4_refclk_clk),                      //   input,    width = 1,       ref_clk_0.clk
		.core_init_n_0   (~rst_controller_reset_out_reset),               //   input,    width = 1,   core_init_n_0.reset_n
		.usr_async_clk_0 (agilex_5_soc_h2f_user1_clk_clk),                //   input,    width = 1, usr_async_clk_0.clk
		.usr_rst_n_0     (emif_bank3a_usr_rst_n_0_reset),                 //  output,    width = 1,     usr_rst_n_0.reset_n
		.s0_axi4_araddr  (mm_interconnect_3_emif_bank3a_s0_axi4_araddr),  //   input,   width = 32,         s0_axi4.araddr
		.s0_axi4_arburst (mm_interconnect_3_emif_bank3a_s0_axi4_arburst), //   input,    width = 2,                .arburst
		.s0_axi4_arid    (mm_interconnect_3_emif_bank3a_s0_axi4_arid),    //   input,    width = 7,                .arid
		.s0_axi4_arlen   (mm_interconnect_3_emif_bank3a_s0_axi4_arlen),   //   input,    width = 8,                .arlen
		.s0_axi4_arlock  (mm_interconnect_3_emif_bank3a_s0_axi4_arlock),  //   input,    width = 1,                .arlock
		.s0_axi4_arqos   (mm_interconnect_3_emif_bank3a_s0_axi4_arqos),   //   input,    width = 4,                .arqos
		.s0_axi4_arsize  (mm_interconnect_3_emif_bank3a_s0_axi4_arsize),  //   input,    width = 3,                .arsize
		.s0_axi4_arvalid (mm_interconnect_3_emif_bank3a_s0_axi4_arvalid), //   input,    width = 1,                .arvalid
		.s0_axi4_aruser  (mm_interconnect_3_emif_bank3a_s0_axi4_aruser),  //   input,   width = 14,                .aruser
		.s0_axi4_arprot  (mm_interconnect_3_emif_bank3a_s0_axi4_arprot),  //   input,    width = 3,                .arprot
		.s0_axi4_awaddr  (mm_interconnect_3_emif_bank3a_s0_axi4_awaddr),  //   input,   width = 32,                .awaddr
		.s0_axi4_awburst (mm_interconnect_3_emif_bank3a_s0_axi4_awburst), //   input,    width = 2,                .awburst
		.s0_axi4_awid    (mm_interconnect_3_emif_bank3a_s0_axi4_awid),    //   input,    width = 7,                .awid
		.s0_axi4_awlen   (mm_interconnect_3_emif_bank3a_s0_axi4_awlen),   //   input,    width = 8,                .awlen
		.s0_axi4_awlock  (mm_interconnect_3_emif_bank3a_s0_axi4_awlock),  //   input,    width = 1,                .awlock
		.s0_axi4_awqos   (mm_interconnect_3_emif_bank3a_s0_axi4_awqos),   //   input,    width = 4,                .awqos
		.s0_axi4_awsize  (mm_interconnect_3_emif_bank3a_s0_axi4_awsize),  //   input,    width = 3,                .awsize
		.s0_axi4_awvalid (mm_interconnect_3_emif_bank3a_s0_axi4_awvalid), //   input,    width = 1,                .awvalid
		.s0_axi4_awuser  (mm_interconnect_3_emif_bank3a_s0_axi4_awuser),  //   input,   width = 14,                .awuser
		.s0_axi4_awprot  (mm_interconnect_3_emif_bank3a_s0_axi4_awprot),  //   input,    width = 3,                .awprot
		.s0_axi4_bready  (mm_interconnect_3_emif_bank3a_s0_axi4_bready),  //   input,    width = 1,                .bready
		.s0_axi4_rready  (mm_interconnect_3_emif_bank3a_s0_axi4_rready),  //   input,    width = 1,                .rready
		.s0_axi4_wdata   (mm_interconnect_3_emif_bank3a_s0_axi4_wdata),   //   input,  width = 256,                .wdata
		.s0_axi4_wstrb   (mm_interconnect_3_emif_bank3a_s0_axi4_wstrb),   //   input,   width = 32,                .wstrb
		.s0_axi4_wlast   (mm_interconnect_3_emif_bank3a_s0_axi4_wlast),   //   input,    width = 1,                .wlast
		.s0_axi4_wvalid  (mm_interconnect_3_emif_bank3a_s0_axi4_wvalid),  //   input,    width = 1,                .wvalid
		.s0_axi4_wuser   (mm_interconnect_3_emif_bank3a_s0_axi4_wuser),   //   input,   width = 64,                .wuser
		.s0_axi4_ruser   (mm_interconnect_3_emif_bank3a_s0_axi4_ruser),   //  output,   width = 64,                .ruser
		.s0_axi4_arready (mm_interconnect_3_emif_bank3a_s0_axi4_arready), //  output,    width = 1,                .arready
		.s0_axi4_awready (mm_interconnect_3_emif_bank3a_s0_axi4_awready), //  output,    width = 1,                .awready
		.s0_axi4_bid     (mm_interconnect_3_emif_bank3a_s0_axi4_bid),     //  output,    width = 7,                .bid
		.s0_axi4_bresp   (mm_interconnect_3_emif_bank3a_s0_axi4_bresp),   //  output,    width = 2,                .bresp
		.s0_axi4_bvalid  (mm_interconnect_3_emif_bank3a_s0_axi4_bvalid),  //  output,    width = 1,                .bvalid
		.s0_axi4_rdata   (mm_interconnect_3_emif_bank3a_s0_axi4_rdata),   //  output,  width = 256,                .rdata
		.s0_axi4_rid     (mm_interconnect_3_emif_bank3a_s0_axi4_rid),     //  output,    width = 7,                .rid
		.s0_axi4_rlast   (mm_interconnect_3_emif_bank3a_s0_axi4_rlast),   //  output,    width = 1,                .rlast
		.s0_axi4_rresp   (mm_interconnect_3_emif_bank3a_s0_axi4_rresp),   //  output,    width = 2,                .rresp
		.s0_axi4_rvalid  (mm_interconnect_3_emif_bank3a_s0_axi4_rvalid),  //  output,    width = 1,                .rvalid
		.s0_axi4_wready  (mm_interconnect_3_emif_bank3a_s0_axi4_wready),  //  output,    width = 1,                .wready
		.mem_ck_t_0      (bank3a_lpddr4_mem_ck_t),                        //  output,    width = 1,           mem_0.mem_ck_t
		.mem_ck_c_0      (bank3a_lpddr4_mem_ck_c),                        //  output,    width = 1,                .mem_ck_c
		.mem_cke_0       (bank3a_lpddr4_mem_cke),                         //  output,    width = 1,                .mem_cke
		.mem_reset_n_0   (bank3a_lpddr4_mem_reset_n),                     //  output,    width = 1,                .mem_reset_n
		.mem_cs_0        (bank3a_lpddr4_mem_cs),                          //  output,    width = 1,                .mem_cs
		.mem_ca_0        (bank3a_lpddr4_mem_ca),                          //  output,    width = 6,                .mem_ca
		.mem_dq_0        (bank3a_lpddr4_mem_dq),                          //   inout,   width = 32,                .mem_dq
		.mem_dqs_t_0     (bank3a_lpddr4_mem_dqs_t),                       //   inout,    width = 4,                .mem_dqs_t
		.mem_dqs_c_0     (bank3a_lpddr4_mem_dqs_c),                       //   inout,    width = 4,                .mem_dqs_c
		.mem_dmi_0       (bank3a_lpddr4_mem_dmi),                         //   inout,    width = 4,                .mem_dmi
		.oct_rzqin_0     (bank3a_lpddr4_oct_oct_rzqin),                   //   input,    width = 1,           oct_0.oct_rzqin
		.s0_axil_clk     (agilex_5_soc_h2f_user1_clk_clk),                //   input,    width = 1,     s0_axil_clk.clk
		.s0_axil_rst_n   (~rst_controller_001_reset_out_reset),           //   input,    width = 1,   s0_axil_rst_n.reset_n
		.s0_axil_awaddr  (mm_interconnect_2_emif_bank3a_s0_axil_awaddr),  //   input,   width = 27,         s0_axil.awaddr
		.s0_axil_awvalid (mm_interconnect_2_emif_bank3a_s0_axil_awvalid), //   input,    width = 1,                .awvalid
		.s0_axil_awready (mm_interconnect_2_emif_bank3a_s0_axil_awready), //  output,    width = 1,                .awready
		.s0_axil_wdata   (mm_interconnect_2_emif_bank3a_s0_axil_wdata),   //   input,   width = 32,                .wdata
		.s0_axil_wstrb   (mm_interconnect_2_emif_bank3a_s0_axil_wstrb),   //   input,    width = 4,                .wstrb
		.s0_axil_wvalid  (mm_interconnect_2_emif_bank3a_s0_axil_wvalid),  //   input,    width = 1,                .wvalid
		.s0_axil_wready  (mm_interconnect_2_emif_bank3a_s0_axil_wready),  //  output,    width = 1,                .wready
		.s0_axil_bresp   (mm_interconnect_2_emif_bank3a_s0_axil_bresp),   //  output,    width = 2,                .bresp
		.s0_axil_bvalid  (mm_interconnect_2_emif_bank3a_s0_axil_bvalid),  //  output,    width = 1,                .bvalid
		.s0_axil_bready  (mm_interconnect_2_emif_bank3a_s0_axil_bready),  //   input,    width = 1,                .bready
		.s0_axil_araddr  (mm_interconnect_2_emif_bank3a_s0_axil_araddr),  //   input,   width = 27,                .araddr
		.s0_axil_arvalid (mm_interconnect_2_emif_bank3a_s0_axil_arvalid), //   input,    width = 1,                .arvalid
		.s0_axil_arready (mm_interconnect_2_emif_bank3a_s0_axil_arready), //  output,    width = 1,                .arready
		.s0_axil_rdata   (mm_interconnect_2_emif_bank3a_s0_axil_rdata),   //  output,   width = 32,                .rdata
		.s0_axil_rresp   (mm_interconnect_2_emif_bank3a_s0_axil_rresp),   //  output,    width = 2,                .rresp
		.s0_axil_rvalid  (mm_interconnect_2_emif_bank3a_s0_axil_rvalid),  //  output,    width = 1,                .rvalid
		.s0_axil_rready  (mm_interconnect_2_emif_bank3a_s0_axil_rready),  //   input,    width = 1,                .rready
		.s0_axil_awprot  (mm_interconnect_2_emif_bank3a_s0_axil_awprot),  //   input,    width = 3,                .awprot
		.s0_axil_arprot  (mm_interconnect_2_emif_bank3a_s0_axil_arprot)   //   input,    width = 3,                .arprot
	);

	ghrd_hps_system_master_2 f2sdram_only_master (
		.clk_clk              (agilex_5_soc_h2f_user1_clk_clk),           //   input,   width = 1,          clk.clk
		.clk_reset_reset      (reset_in_out_reset_reset),                 //   input,   width = 1,    clk_reset.reset
		.master_reset_reset   (),                                         //  output,   width = 1, master_reset.reset
		.master_address       (f2sdram_only_master_master_address),       //  output,  width = 32,       master.address
		.master_readdata      (f2sdram_only_master_master_readdata),      //   input,  width = 32,             .readdata
		.master_read          (f2sdram_only_master_master_read),          //  output,   width = 1,             .read
		.master_write         (f2sdram_only_master_master_write),         //  output,   width = 1,             .write
		.master_writedata     (f2sdram_only_master_master_writedata),     //  output,  width = 32,             .writedata
		.master_waitrequest   (f2sdram_only_master_master_waitrequest),   //   input,   width = 1,             .waitrequest
		.master_readdatavalid (f2sdram_only_master_master_readdatavalid), //   input,   width = 1,             .readdatavalid
		.master_byteenable    (f2sdram_only_master_master_byteenable)     //  output,   width = 4,             .byteenable
	);

	ghrd_hps_system_master_1 fpga_only_master (
		.clk_clk              (agilex_5_soc_h2f_user1_clk_clk),        //   input,   width = 1,          clk.clk
		.clk_reset_reset      (rst_controller_002_reset_out_reset),    //   input,   width = 1,    clk_reset.reset
		.master_reset_reset   (fpga_only_master_master_reset_reset),   //  output,   width = 1, master_reset.reset
		.master_address       (fpga_only_master_master_address),       //  output,  width = 32,       master.address
		.master_readdata      (fpga_only_master_master_readdata),      //   input,  width = 32,             .readdata
		.master_read          (fpga_only_master_master_read),          //  output,   width = 1,             .read
		.master_write         (fpga_only_master_master_write),         //  output,   width = 1,             .write
		.master_writedata     (fpga_only_master_master_writedata),     //  output,  width = 32,             .writedata
		.master_waitrequest   (fpga_only_master_master_waitrequest),   //   input,   width = 1,             .waitrequest
		.master_readdatavalid (fpga_only_master_master_readdatavalid), //   input,   width = 1,             .readdatavalid
		.master_byteenable    (fpga_only_master_master_byteenable)     //  output,   width = 4,             .byteenable
	);

	ghrd_hps_system_intel_onchip_memory_0 onchip_sram (
		.clk        (agilex_5_soc_h2f_user0_clk_clk),               //   input,   width = 1,   clk1.clk
		.s1_arid    (mm_interconnect_1_onchip_sram_axi_s1_arid),    //   input,   width = 7, axi_s1.arid
		.s1_araddr  (mm_interconnect_1_onchip_sram_axi_s1_araddr),  //   input,  width = 15,       .araddr
		.s1_arlen   (mm_interconnect_1_onchip_sram_axi_s1_arlen),   //   input,   width = 8,       .arlen
		.s1_arsize  (mm_interconnect_1_onchip_sram_axi_s1_arsize),  //   input,   width = 3,       .arsize
		.s1_arburst (mm_interconnect_1_onchip_sram_axi_s1_arburst), //   input,   width = 2,       .arburst
		.s1_arready (mm_interconnect_1_onchip_sram_axi_s1_arready), //  output,   width = 1,       .arready
		.s1_arvalid (mm_interconnect_1_onchip_sram_axi_s1_arvalid), //   input,   width = 1,       .arvalid
		.s1_awid    (mm_interconnect_1_onchip_sram_axi_s1_awid),    //   input,   width = 7,       .awid
		.s1_awaddr  (mm_interconnect_1_onchip_sram_axi_s1_awaddr),  //   input,  width = 15,       .awaddr
		.s1_awlen   (mm_interconnect_1_onchip_sram_axi_s1_awlen),   //   input,   width = 8,       .awlen
		.s1_awsize  (mm_interconnect_1_onchip_sram_axi_s1_awsize),  //   input,   width = 3,       .awsize
		.s1_awburst (mm_interconnect_1_onchip_sram_axi_s1_awburst), //   input,   width = 2,       .awburst
		.s1_awready (mm_interconnect_1_onchip_sram_axi_s1_awready), //  output,   width = 1,       .awready
		.s1_awvalid (mm_interconnect_1_onchip_sram_axi_s1_awvalid), //   input,   width = 1,       .awvalid
		.s1_rid     (mm_interconnect_1_onchip_sram_axi_s1_rid),     //  output,   width = 7,       .rid
		.s1_rdata   (mm_interconnect_1_onchip_sram_axi_s1_rdata),   //  output,  width = 64,       .rdata
		.s1_rlast   (mm_interconnect_1_onchip_sram_axi_s1_rlast),   //  output,   width = 1,       .rlast
		.s1_rready  (mm_interconnect_1_onchip_sram_axi_s1_rready),  //   input,   width = 1,       .rready
		.s1_rvalid  (mm_interconnect_1_onchip_sram_axi_s1_rvalid),  //  output,   width = 1,       .rvalid
		.s1_rresp   (mm_interconnect_1_onchip_sram_axi_s1_rresp),   //  output,   width = 2,       .rresp
		.s1_wdata   (mm_interconnect_1_onchip_sram_axi_s1_wdata),   //   input,  width = 64,       .wdata
		.s1_wstrb   (mm_interconnect_1_onchip_sram_axi_s1_wstrb),   //   input,   width = 8,       .wstrb
		.s1_wlast   (mm_interconnect_1_onchip_sram_axi_s1_wlast),   //   input,   width = 1,       .wlast
		.s1_wready  (mm_interconnect_1_onchip_sram_axi_s1_wready),  //  output,   width = 1,       .wready
		.s1_wvalid  (mm_interconnect_1_onchip_sram_axi_s1_wvalid),  //   input,   width = 1,       .wvalid
		.s1_bid     (mm_interconnect_1_onchip_sram_axi_s1_bid),     //  output,   width = 7,       .bid
		.s1_bresp   (mm_interconnect_1_onchip_sram_axi_s1_bresp),   //  output,   width = 2,       .bresp
		.s1_bready  (mm_interconnect_1_onchip_sram_axi_s1_bready),  //   input,   width = 1,       .bready
		.s1_bvalid  (mm_interconnect_1_onchip_sram_axi_s1_bvalid),  //  output,   width = 1,       .bvalid
		.reset      (rst_controller_003_reset_out_reset)            //   input,   width = 1, reset1.reset
	);

	ghrd_hps_system_reset_in reset_in (
		.clk       (agilex_5_soc_h2f_user1_clk_clk), //   input,  width = 1,       clk.clk
		.in_reset  (sys_reset_reset),                //   input,  width = 1,  in_reset.reset
		.out_reset (reset_in_out_reset_reset)        //  output,  width = 1, out_reset.reset
	);

	peripheral_sys peripheral_sys_0 (
		.clk_clk                               (agilex_5_soc_h2f_user1_clk_clk),                                           //   input,   width = 1,                     clk.clk
		.dipsw_export                          (dipsw_export),                                                             //   input,   width = 2,                   dipsw.export
		.dipsw_irq_irq                         (irq_mapper_receiver0_irq),                                                 //  output,   width = 1,               dipsw_irq.irq
		.jtag_uart_irq_irq                     (irq_mapper_receiver2_irq),                                                 //  output,   width = 1,           jtag_uart_irq.irq
		.mm_peripheral_bridge_s0_waitrequest   (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_waitrequest),   //  output,   width = 1, mm_peripheral_bridge_s0.waitrequest
		.mm_peripheral_bridge_s0_readdata      (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_readdata),      //  output,  width = 32,                        .readdata
		.mm_peripheral_bridge_s0_readdatavalid (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_readdatavalid), //  output,   width = 1,                        .readdatavalid
		.mm_peripheral_bridge_s0_burstcount    (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_burstcount),    //   input,   width = 1,                        .burstcount
		.mm_peripheral_bridge_s0_writedata     (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_writedata),     //   input,  width = 32,                        .writedata
		.mm_peripheral_bridge_s0_address       (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_address),       //   input,  width = 24,                        .address
		.mm_peripheral_bridge_s0_write         (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_write),         //   input,   width = 1,                        .write
		.mm_peripheral_bridge_s0_read          (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_read),          //   input,   width = 1,                        .read
		.mm_peripheral_bridge_s0_byteenable    (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_byteenable),    //   input,   width = 4,                        .byteenable
		.mm_peripheral_bridge_s0_debugaccess   (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_debugaccess),   //   input,   width = 1,                        .debugaccess
		.pb_export                             (pb_export),                                                                //   input,   width = 2,                      pb.export
		.pb_irq_irq                            (irq_mapper_receiver3_irq),                                                 //  output,   width = 1,                  pb_irq.irq
		.reset_reset                           (reset_in_out_reset_reset),                                                 //   input,   width = 1,                   reset.reset
		.rgb_led0_export                       (rgb_led0_export),                                                          //  output,   width = 3,                rgb_led0.export
		.rgb_led1_export                       (rgb_led1_export),                                                          //  output,   width = 3,                rgb_led1.export
		.rgb_led2_export                       (rgb_led2_export),                                                          //  output,   width = 3,                rgb_led2.export
		.rgb_led3_export                       (rgb_led3_export)                                                           //  output,   width = 3,                rgb_led3.export
	);

	video_sys video_sys_0 (
		.hdmi_h_clk                       (hdmi_h_clk),                                                     //  output,   width = 1,               hdmi.h_clk
		.hdmi_h16_hsync                   (hdmi_h16_hsync),                                                 //  output,   width = 1,                   .h16_hsync
		.hdmi_h16_vsync                   (hdmi_h16_vsync),                                                 //  output,   width = 1,                   .h16_vsync
		.hdmi_h16_data_e                  (hdmi_h16_data_e),                                                //  output,   width = 1,                   .h16_data_e
		.hdmi_h16_data                    (hdmi_h16_data),                                                  //  output,  width = 16,                   .h16_data
		.hdmi_h16_es_data                 (hdmi_h16_es_data),                                               //  output,  width = 16,                   .h16_es_data
		.hdmi_h24_hsync                   (hdmi_h24_hsync),                                                 //  output,   width = 1,                   .h24_hsync
		.hdmi_h24_vsync                   (hdmi_h24_vsync),                                                 //  output,   width = 1,                   .h24_vsync
		.hdmi_h24_data_e                  (hdmi_h24_data_e),                                                //  output,   width = 1,                   .h24_data_e
		.hdmi_h24_data                    (hdmi_h24_data),                                                  //  output,  width = 24,                   .h24_data
		.hdmi_h36_hsync                   (hdmi_h36_hsync),                                                 //  output,   width = 1,                   .h36_hsync
		.hdmi_h36_vsync                   (hdmi_h36_vsync),                                                 //  output,   width = 1,                   .h36_vsync
		.hdmi_h36_data_e                  (hdmi_h36_data_e),                                                //  output,   width = 1,                   .h36_data_e
		.hdmi_h36_data                    (hdmi_h36_data),                                                  //  output,  width = 36,                   .h36_data
		.clk_clk                          (agilex_5_soc_h2f_user1_clk_clk),                                 //   input,   width = 1,                clk.clk
		.hdmi_dmac_irq                    (irq_mapper_receiver1_irq),                                       //  output,   width = 1,          hdmi_dmac.irq
		.hdmi_dmac_master_awvalid         (video_sys_0_hdmi_dmac_master_awvalid),                           //  output,   width = 1,   hdmi_dmac_master.awvalid
		.hdmi_dmac_master_awaddr          (video_sys_0_hdmi_dmac_master_awaddr),                            //  output,  width = 32,                   .awaddr
		.hdmi_dmac_master_awready         (video_sys_0_hdmi_dmac_master_awready),                           //   input,   width = 1,                   .awready
		.hdmi_dmac_master_wvalid          (video_sys_0_hdmi_dmac_master_wvalid),                            //  output,   width = 1,                   .wvalid
		.hdmi_dmac_master_wdata           (video_sys_0_hdmi_dmac_master_wdata),                             //  output,  width = 64,                   .wdata
		.hdmi_dmac_master_wstrb           (video_sys_0_hdmi_dmac_master_wstrb),                             //  output,   width = 8,                   .wstrb
		.hdmi_dmac_master_wready          (video_sys_0_hdmi_dmac_master_wready),                            //   input,   width = 1,                   .wready
		.hdmi_dmac_master_bvalid          (video_sys_0_hdmi_dmac_master_bvalid),                            //   input,   width = 1,                   .bvalid
		.hdmi_dmac_master_bresp           (video_sys_0_hdmi_dmac_master_bresp),                             //   input,   width = 2,                   .bresp
		.hdmi_dmac_master_bready          (video_sys_0_hdmi_dmac_master_bready),                            //  output,   width = 1,                   .bready
		.hdmi_dmac_master_arvalid         (video_sys_0_hdmi_dmac_master_arvalid),                           //  output,   width = 1,                   .arvalid
		.hdmi_dmac_master_araddr          (video_sys_0_hdmi_dmac_master_araddr),                            //  output,  width = 32,                   .araddr
		.hdmi_dmac_master_arready         (video_sys_0_hdmi_dmac_master_arready),                           //   input,   width = 1,                   .arready
		.hdmi_dmac_master_rvalid          (video_sys_0_hdmi_dmac_master_rvalid),                            //   input,   width = 1,                   .rvalid
		.hdmi_dmac_master_rresp           (video_sys_0_hdmi_dmac_master_rresp),                             //   input,   width = 2,                   .rresp
		.hdmi_dmac_master_rdata           (video_sys_0_hdmi_dmac_master_rdata),                             //   input,  width = 64,                   .rdata
		.hdmi_dmac_master_rready          (video_sys_0_hdmi_dmac_master_rready),                            //  output,   width = 1,                   .rready
		.hdmi_dmac_master_awlen           (video_sys_0_hdmi_dmac_master_awlen),                             //  output,   width = 4,                   .awlen
		.hdmi_dmac_master_awsize          (video_sys_0_hdmi_dmac_master_awsize),                            //  output,   width = 3,                   .awsize
		.hdmi_dmac_master_awburst         (video_sys_0_hdmi_dmac_master_awburst),                           //  output,   width = 2,                   .awburst
		.hdmi_dmac_master_awcache         (video_sys_0_hdmi_dmac_master_awcache),                           //  output,   width = 4,                   .awcache
		.hdmi_dmac_master_awprot          (video_sys_0_hdmi_dmac_master_awprot),                            //  output,   width = 3,                   .awprot
		.hdmi_dmac_master_wlast           (video_sys_0_hdmi_dmac_master_wlast),                             //  output,   width = 1,                   .wlast
		.hdmi_dmac_master_arlen           (video_sys_0_hdmi_dmac_master_arlen),                             //  output,   width = 4,                   .arlen
		.hdmi_dmac_master_arsize          (video_sys_0_hdmi_dmac_master_arsize),                            //  output,   width = 3,                   .arsize
		.hdmi_dmac_master_arburst         (video_sys_0_hdmi_dmac_master_arburst),                           //  output,   width = 2,                   .arburst
		.hdmi_dmac_master_arcache         (video_sys_0_hdmi_dmac_master_arcache),                           //  output,   width = 4,                   .arcache
		.hdmi_dmac_master_arprot          (video_sys_0_hdmi_dmac_master_arprot),                            //  output,   width = 3,                   .arprot
		.hdmi_dmac_master_awid            (video_sys_0_hdmi_dmac_master_awid),                              //  output,   width = 1,                   .awid
		.hdmi_dmac_master_awlock          (video_sys_0_hdmi_dmac_master_awlock),                            //  output,   width = 2,                   .awlock
		.hdmi_dmac_master_wid             (video_sys_0_hdmi_dmac_master_wid),                               //  output,   width = 1,                   .wid
		.hdmi_dmac_master_arid            (video_sys_0_hdmi_dmac_master_arid),                              //  output,   width = 1,                   .arid
		.hdmi_dmac_master_arlock          (video_sys_0_hdmi_dmac_master_arlock),                            //  output,   width = 2,                   .arlock
		.hdmi_dmac_master_rid             (video_sys_0_hdmi_dmac_master_rid),                               //   input,   width = 1,                   .rid
		.hdmi_dmac_master_bid             (video_sys_0_hdmi_dmac_master_bid),                               //   input,   width = 1,                   .bid
		.hdmi_dmac_master_rlast           (video_sys_0_hdmi_dmac_master_rlast),                             //   input,   width = 1,                   .rlast
		.hdmi_pll_refclk_clk              (hdmi_pll_refclk_clk),                                            //   input,   width = 1,    hdmi_pll_refclk.clk
		.mm_video_bridge_s0_waitrequest   (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_waitrequest),   //  output,   width = 1, mm_video_bridge_s0.waitrequest
		.mm_video_bridge_s0_readdata      (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_readdata),      //  output,  width = 32,                   .readdata
		.mm_video_bridge_s0_readdatavalid (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_readdatavalid), //  output,   width = 1,                   .readdatavalid
		.mm_video_bridge_s0_burstcount    (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_burstcount),    //   input,   width = 1,                   .burstcount
		.mm_video_bridge_s0_writedata     (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_writedata),     //   input,  width = 32,                   .writedata
		.mm_video_bridge_s0_address       (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_address),       //   input,  width = 24,                   .address
		.mm_video_bridge_s0_write         (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_write),         //   input,   width = 1,                   .write
		.mm_video_bridge_s0_read          (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_read),          //   input,   width = 1,                   .read
		.mm_video_bridge_s0_byteenable    (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_byteenable),    //   input,   width = 4,                   .byteenable
		.mm_video_bridge_s0_debugaccess   (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_debugaccess),   //   input,   width = 1,                   .debugaccess
		.reset_reset                      (reset_in_out_reset_reset)                                        //   input,   width = 1,              reset.reset
	);

	ghrd_hps_system_altera_mm_interconnect_1920_52h6z3a mm_interconnect_0 (
		.f2sdram_only_master_master_address                                      (f2sdram_only_master_master_address),              //   input,  width = 32,                                        f2sdram_only_master_master.address
		.f2sdram_only_master_master_waitrequest                                  (f2sdram_only_master_master_waitrequest),          //  output,   width = 1,                                                                  .waitrequest
		.f2sdram_only_master_master_byteenable                                   (f2sdram_only_master_master_byteenable),           //   input,   width = 4,                                                                  .byteenable
		.f2sdram_only_master_master_read                                         (f2sdram_only_master_master_read),                 //   input,   width = 1,                                                                  .read
		.f2sdram_only_master_master_readdata                                     (f2sdram_only_master_master_readdata),             //  output,  width = 32,                                                                  .readdata
		.f2sdram_only_master_master_readdatavalid                                (f2sdram_only_master_master_readdatavalid),        //  output,   width = 1,                                                                  .readdatavalid
		.f2sdram_only_master_master_write                                        (f2sdram_only_master_master_write),                //   input,   width = 1,                                                                  .write
		.f2sdram_only_master_master_writedata                                    (f2sdram_only_master_master_writedata),            //   input,  width = 32,                                                                  .writedata
		.agilex_5_soc_f2sdram_awid                                               (mm_interconnect_0_agilex_5_soc_f2sdram_awid),     //  output,   width = 5,                                              agilex_5_soc_f2sdram.awid
		.agilex_5_soc_f2sdram_awaddr                                             (mm_interconnect_0_agilex_5_soc_f2sdram_awaddr),   //  output,  width = 32,                                                                  .awaddr
		.agilex_5_soc_f2sdram_awlen                                              (mm_interconnect_0_agilex_5_soc_f2sdram_awlen),    //  output,   width = 8,                                                                  .awlen
		.agilex_5_soc_f2sdram_awsize                                             (mm_interconnect_0_agilex_5_soc_f2sdram_awsize),   //  output,   width = 3,                                                                  .awsize
		.agilex_5_soc_f2sdram_awburst                                            (mm_interconnect_0_agilex_5_soc_f2sdram_awburst),  //  output,   width = 2,                                                                  .awburst
		.agilex_5_soc_f2sdram_awlock                                             (mm_interconnect_0_agilex_5_soc_f2sdram_awlock),   //  output,   width = 1,                                                                  .awlock
		.agilex_5_soc_f2sdram_awcache                                            (mm_interconnect_0_agilex_5_soc_f2sdram_awcache),  //  output,   width = 4,                                                                  .awcache
		.agilex_5_soc_f2sdram_awprot                                             (mm_interconnect_0_agilex_5_soc_f2sdram_awprot),   //  output,   width = 3,                                                                  .awprot
		.agilex_5_soc_f2sdram_awuser                                             (mm_interconnect_0_agilex_5_soc_f2sdram_awuser),   //  output,   width = 8,                                                                  .awuser
		.agilex_5_soc_f2sdram_awqos                                              (mm_interconnect_0_agilex_5_soc_f2sdram_awqos),    //  output,   width = 4,                                                                  .awqos
		.agilex_5_soc_f2sdram_awregion                                           (mm_interconnect_0_agilex_5_soc_f2sdram_awregion), //  output,   width = 4,                                                                  .awregion
		.agilex_5_soc_f2sdram_awvalid                                            (mm_interconnect_0_agilex_5_soc_f2sdram_awvalid),  //  output,   width = 1,                                                                  .awvalid
		.agilex_5_soc_f2sdram_awready                                            (mm_interconnect_0_agilex_5_soc_f2sdram_awready),  //   input,   width = 1,                                                                  .awready
		.agilex_5_soc_f2sdram_wdata                                              (mm_interconnect_0_agilex_5_soc_f2sdram_wdata),    //  output,  width = 64,                                                                  .wdata
		.agilex_5_soc_f2sdram_wstrb                                              (mm_interconnect_0_agilex_5_soc_f2sdram_wstrb),    //  output,   width = 8,                                                                  .wstrb
		.agilex_5_soc_f2sdram_wlast                                              (mm_interconnect_0_agilex_5_soc_f2sdram_wlast),    //  output,   width = 1,                                                                  .wlast
		.agilex_5_soc_f2sdram_wvalid                                             (mm_interconnect_0_agilex_5_soc_f2sdram_wvalid),   //  output,   width = 1,                                                                  .wvalid
		.agilex_5_soc_f2sdram_wuser                                              (mm_interconnect_0_agilex_5_soc_f2sdram_wuser),    //  output,   width = 8,                                                                  .wuser
		.agilex_5_soc_f2sdram_wready                                             (mm_interconnect_0_agilex_5_soc_f2sdram_wready),   //   input,   width = 1,                                                                  .wready
		.agilex_5_soc_f2sdram_bid                                                (mm_interconnect_0_agilex_5_soc_f2sdram_bid),      //   input,   width = 5,                                                                  .bid
		.agilex_5_soc_f2sdram_bresp                                              (mm_interconnect_0_agilex_5_soc_f2sdram_bresp),    //   input,   width = 2,                                                                  .bresp
		.agilex_5_soc_f2sdram_buser                                              (mm_interconnect_0_agilex_5_soc_f2sdram_buser),    //   input,   width = 8,                                                                  .buser
		.agilex_5_soc_f2sdram_bvalid                                             (mm_interconnect_0_agilex_5_soc_f2sdram_bvalid),   //   input,   width = 1,                                                                  .bvalid
		.agilex_5_soc_f2sdram_bready                                             (mm_interconnect_0_agilex_5_soc_f2sdram_bready),   //  output,   width = 1,                                                                  .bready
		.agilex_5_soc_f2sdram_arid                                               (mm_interconnect_0_agilex_5_soc_f2sdram_arid),     //  output,   width = 5,                                                                  .arid
		.agilex_5_soc_f2sdram_araddr                                             (mm_interconnect_0_agilex_5_soc_f2sdram_araddr),   //  output,  width = 32,                                                                  .araddr
		.agilex_5_soc_f2sdram_arlen                                              (mm_interconnect_0_agilex_5_soc_f2sdram_arlen),    //  output,   width = 8,                                                                  .arlen
		.agilex_5_soc_f2sdram_arsize                                             (mm_interconnect_0_agilex_5_soc_f2sdram_arsize),   //  output,   width = 3,                                                                  .arsize
		.agilex_5_soc_f2sdram_arburst                                            (mm_interconnect_0_agilex_5_soc_f2sdram_arburst),  //  output,   width = 2,                                                                  .arburst
		.agilex_5_soc_f2sdram_arlock                                             (mm_interconnect_0_agilex_5_soc_f2sdram_arlock),   //  output,   width = 1,                                                                  .arlock
		.agilex_5_soc_f2sdram_arcache                                            (mm_interconnect_0_agilex_5_soc_f2sdram_arcache),  //  output,   width = 4,                                                                  .arcache
		.agilex_5_soc_f2sdram_arprot                                             (mm_interconnect_0_agilex_5_soc_f2sdram_arprot),   //  output,   width = 3,                                                                  .arprot
		.agilex_5_soc_f2sdram_aruser                                             (mm_interconnect_0_agilex_5_soc_f2sdram_aruser),   //  output,   width = 8,                                                                  .aruser
		.agilex_5_soc_f2sdram_arqos                                              (mm_interconnect_0_agilex_5_soc_f2sdram_arqos),    //  output,   width = 4,                                                                  .arqos
		.agilex_5_soc_f2sdram_arregion                                           (mm_interconnect_0_agilex_5_soc_f2sdram_arregion), //  output,   width = 4,                                                                  .arregion
		.agilex_5_soc_f2sdram_arvalid                                            (mm_interconnect_0_agilex_5_soc_f2sdram_arvalid),  //  output,   width = 1,                                                                  .arvalid
		.agilex_5_soc_f2sdram_arready                                            (mm_interconnect_0_agilex_5_soc_f2sdram_arready),  //   input,   width = 1,                                                                  .arready
		.agilex_5_soc_f2sdram_rid                                                (mm_interconnect_0_agilex_5_soc_f2sdram_rid),      //   input,   width = 5,                                                                  .rid
		.agilex_5_soc_f2sdram_rdata                                              (mm_interconnect_0_agilex_5_soc_f2sdram_rdata),    //   input,  width = 64,                                                                  .rdata
		.agilex_5_soc_f2sdram_rresp                                              (mm_interconnect_0_agilex_5_soc_f2sdram_rresp),    //   input,   width = 2,                                                                  .rresp
		.agilex_5_soc_f2sdram_rlast                                              (mm_interconnect_0_agilex_5_soc_f2sdram_rlast),    //   input,   width = 1,                                                                  .rlast
		.agilex_5_soc_f2sdram_rvalid                                             (mm_interconnect_0_agilex_5_soc_f2sdram_rvalid),   //   input,   width = 1,                                                                  .rvalid
		.agilex_5_soc_f2sdram_rready                                             (mm_interconnect_0_agilex_5_soc_f2sdram_rready),   //  output,   width = 1,                                                                  .rready
		.agilex_5_soc_f2sdram_ruser                                              (mm_interconnect_0_agilex_5_soc_f2sdram_ruser),    //   input,   width = 8,                                                                  .ruser
		.video_sys_0_hdmi_dmac_master_awid                                       (video_sys_0_hdmi_dmac_master_awid),               //   input,   width = 1,                                      video_sys_0_hdmi_dmac_master.awid
		.video_sys_0_hdmi_dmac_master_awaddr                                     (video_sys_0_hdmi_dmac_master_awaddr),             //   input,  width = 32,                                                                  .awaddr
		.video_sys_0_hdmi_dmac_master_awlen                                      (video_sys_0_hdmi_dmac_master_awlen),              //   input,   width = 4,                                                                  .awlen
		.video_sys_0_hdmi_dmac_master_awsize                                     (video_sys_0_hdmi_dmac_master_awsize),             //   input,   width = 3,                                                                  .awsize
		.video_sys_0_hdmi_dmac_master_awburst                                    (video_sys_0_hdmi_dmac_master_awburst),            //   input,   width = 2,                                                                  .awburst
		.video_sys_0_hdmi_dmac_master_awlock                                     (video_sys_0_hdmi_dmac_master_awlock),             //   input,   width = 2,                                                                  .awlock
		.video_sys_0_hdmi_dmac_master_awcache                                    (video_sys_0_hdmi_dmac_master_awcache),            //   input,   width = 4,                                                                  .awcache
		.video_sys_0_hdmi_dmac_master_awprot                                     (video_sys_0_hdmi_dmac_master_awprot),             //   input,   width = 3,                                                                  .awprot
		.video_sys_0_hdmi_dmac_master_awvalid                                    (video_sys_0_hdmi_dmac_master_awvalid),            //   input,   width = 1,                                                                  .awvalid
		.video_sys_0_hdmi_dmac_master_awready                                    (video_sys_0_hdmi_dmac_master_awready),            //  output,   width = 1,                                                                  .awready
		.video_sys_0_hdmi_dmac_master_wid                                        (video_sys_0_hdmi_dmac_master_wid),                //   input,   width = 1,                                                                  .wid
		.video_sys_0_hdmi_dmac_master_wdata                                      (video_sys_0_hdmi_dmac_master_wdata),              //   input,  width = 64,                                                                  .wdata
		.video_sys_0_hdmi_dmac_master_wstrb                                      (video_sys_0_hdmi_dmac_master_wstrb),              //   input,   width = 8,                                                                  .wstrb
		.video_sys_0_hdmi_dmac_master_wlast                                      (video_sys_0_hdmi_dmac_master_wlast),              //   input,   width = 1,                                                                  .wlast
		.video_sys_0_hdmi_dmac_master_wvalid                                     (video_sys_0_hdmi_dmac_master_wvalid),             //   input,   width = 1,                                                                  .wvalid
		.video_sys_0_hdmi_dmac_master_wready                                     (video_sys_0_hdmi_dmac_master_wready),             //  output,   width = 1,                                                                  .wready
		.video_sys_0_hdmi_dmac_master_bid                                        (video_sys_0_hdmi_dmac_master_bid),                //  output,   width = 1,                                                                  .bid
		.video_sys_0_hdmi_dmac_master_bresp                                      (video_sys_0_hdmi_dmac_master_bresp),              //  output,   width = 2,                                                                  .bresp
		.video_sys_0_hdmi_dmac_master_bvalid                                     (video_sys_0_hdmi_dmac_master_bvalid),             //  output,   width = 1,                                                                  .bvalid
		.video_sys_0_hdmi_dmac_master_bready                                     (video_sys_0_hdmi_dmac_master_bready),             //   input,   width = 1,                                                                  .bready
		.video_sys_0_hdmi_dmac_master_arid                                       (video_sys_0_hdmi_dmac_master_arid),               //   input,   width = 1,                                                                  .arid
		.video_sys_0_hdmi_dmac_master_araddr                                     (video_sys_0_hdmi_dmac_master_araddr),             //   input,  width = 32,                                                                  .araddr
		.video_sys_0_hdmi_dmac_master_arlen                                      (video_sys_0_hdmi_dmac_master_arlen),              //   input,   width = 4,                                                                  .arlen
		.video_sys_0_hdmi_dmac_master_arsize                                     (video_sys_0_hdmi_dmac_master_arsize),             //   input,   width = 3,                                                                  .arsize
		.video_sys_0_hdmi_dmac_master_arburst                                    (video_sys_0_hdmi_dmac_master_arburst),            //   input,   width = 2,                                                                  .arburst
		.video_sys_0_hdmi_dmac_master_arlock                                     (video_sys_0_hdmi_dmac_master_arlock),             //   input,   width = 2,                                                                  .arlock
		.video_sys_0_hdmi_dmac_master_arcache                                    (video_sys_0_hdmi_dmac_master_arcache),            //   input,   width = 4,                                                                  .arcache
		.video_sys_0_hdmi_dmac_master_arprot                                     (video_sys_0_hdmi_dmac_master_arprot),             //   input,   width = 3,                                                                  .arprot
		.video_sys_0_hdmi_dmac_master_arvalid                                    (video_sys_0_hdmi_dmac_master_arvalid),            //   input,   width = 1,                                                                  .arvalid
		.video_sys_0_hdmi_dmac_master_arready                                    (video_sys_0_hdmi_dmac_master_arready),            //  output,   width = 1,                                                                  .arready
		.video_sys_0_hdmi_dmac_master_rid                                        (video_sys_0_hdmi_dmac_master_rid),                //  output,   width = 1,                                                                  .rid
		.video_sys_0_hdmi_dmac_master_rdata                                      (video_sys_0_hdmi_dmac_master_rdata),              //  output,  width = 64,                                                                  .rdata
		.video_sys_0_hdmi_dmac_master_rresp                                      (video_sys_0_hdmi_dmac_master_rresp),              //  output,   width = 2,                                                                  .rresp
		.video_sys_0_hdmi_dmac_master_rlast                                      (video_sys_0_hdmi_dmac_master_rlast),              //  output,   width = 1,                                                                  .rlast
		.video_sys_0_hdmi_dmac_master_rvalid                                     (video_sys_0_hdmi_dmac_master_rvalid),             //  output,   width = 1,                                                                  .rvalid
		.video_sys_0_hdmi_dmac_master_rready                                     (video_sys_0_hdmi_dmac_master_rready),             //   input,   width = 1,                                                                  .rready
		.f2sdram_only_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),              //   input,   width = 1, f2sdram_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.agilex_5_soc_h2f_user1_clk_clk                                          (agilex_5_soc_h2f_user1_clk_clk)                   //   input,   width = 1,                                        agilex_5_soc_h2f_user1_clk.clk
	);

	ghrd_hps_system_altera_mm_interconnect_1920_ei2j4cq mm_interconnect_1 (
		.agilex_5_soc_hps2fpga_awid                                             (agilex_5_soc_hps2fpga_awid),                                               //   input,   width = 4,                                            agilex_5_soc_hps2fpga.awid
		.agilex_5_soc_hps2fpga_awaddr                                           (agilex_5_soc_hps2fpga_awaddr),                                             //   input,  width = 32,                                                                 .awaddr
		.agilex_5_soc_hps2fpga_awlen                                            (agilex_5_soc_hps2fpga_awlen),                                              //   input,   width = 8,                                                                 .awlen
		.agilex_5_soc_hps2fpga_awsize                                           (agilex_5_soc_hps2fpga_awsize),                                             //   input,   width = 3,                                                                 .awsize
		.agilex_5_soc_hps2fpga_awburst                                          (agilex_5_soc_hps2fpga_awburst),                                            //   input,   width = 2,                                                                 .awburst
		.agilex_5_soc_hps2fpga_awlock                                           (agilex_5_soc_hps2fpga_awlock),                                             //   input,   width = 1,                                                                 .awlock
		.agilex_5_soc_hps2fpga_awcache                                          (agilex_5_soc_hps2fpga_awcache),                                            //   input,   width = 4,                                                                 .awcache
		.agilex_5_soc_hps2fpga_awprot                                           (agilex_5_soc_hps2fpga_awprot),                                             //   input,   width = 3,                                                                 .awprot
		.agilex_5_soc_hps2fpga_awvalid                                          (agilex_5_soc_hps2fpga_awvalid),                                            //   input,   width = 1,                                                                 .awvalid
		.agilex_5_soc_hps2fpga_awready                                          (agilex_5_soc_hps2fpga_awready),                                            //  output,   width = 1,                                                                 .awready
		.agilex_5_soc_hps2fpga_wdata                                            (agilex_5_soc_hps2fpga_wdata),                                              //   input,  width = 32,                                                                 .wdata
		.agilex_5_soc_hps2fpga_wstrb                                            (agilex_5_soc_hps2fpga_wstrb),                                              //   input,   width = 4,                                                                 .wstrb
		.agilex_5_soc_hps2fpga_wlast                                            (agilex_5_soc_hps2fpga_wlast),                                              //   input,   width = 1,                                                                 .wlast
		.agilex_5_soc_hps2fpga_wvalid                                           (agilex_5_soc_hps2fpga_wvalid),                                             //   input,   width = 1,                                                                 .wvalid
		.agilex_5_soc_hps2fpga_wready                                           (agilex_5_soc_hps2fpga_wready),                                             //  output,   width = 1,                                                                 .wready
		.agilex_5_soc_hps2fpga_bid                                              (agilex_5_soc_hps2fpga_bid),                                                //  output,   width = 4,                                                                 .bid
		.agilex_5_soc_hps2fpga_bresp                                            (agilex_5_soc_hps2fpga_bresp),                                              //  output,   width = 2,                                                                 .bresp
		.agilex_5_soc_hps2fpga_bvalid                                           (agilex_5_soc_hps2fpga_bvalid),                                             //  output,   width = 1,                                                                 .bvalid
		.agilex_5_soc_hps2fpga_bready                                           (agilex_5_soc_hps2fpga_bready),                                             //   input,   width = 1,                                                                 .bready
		.agilex_5_soc_hps2fpga_arid                                             (agilex_5_soc_hps2fpga_arid),                                               //   input,   width = 4,                                                                 .arid
		.agilex_5_soc_hps2fpga_araddr                                           (agilex_5_soc_hps2fpga_araddr),                                             //   input,  width = 32,                                                                 .araddr
		.agilex_5_soc_hps2fpga_arlen                                            (agilex_5_soc_hps2fpga_arlen),                                              //   input,   width = 8,                                                                 .arlen
		.agilex_5_soc_hps2fpga_arsize                                           (agilex_5_soc_hps2fpga_arsize),                                             //   input,   width = 3,                                                                 .arsize
		.agilex_5_soc_hps2fpga_arburst                                          (agilex_5_soc_hps2fpga_arburst),                                            //   input,   width = 2,                                                                 .arburst
		.agilex_5_soc_hps2fpga_arlock                                           (agilex_5_soc_hps2fpga_arlock),                                             //   input,   width = 1,                                                                 .arlock
		.agilex_5_soc_hps2fpga_arcache                                          (agilex_5_soc_hps2fpga_arcache),                                            //   input,   width = 4,                                                                 .arcache
		.agilex_5_soc_hps2fpga_arprot                                           (agilex_5_soc_hps2fpga_arprot),                                             //   input,   width = 3,                                                                 .arprot
		.agilex_5_soc_hps2fpga_arvalid                                          (agilex_5_soc_hps2fpga_arvalid),                                            //   input,   width = 1,                                                                 .arvalid
		.agilex_5_soc_hps2fpga_arready                                          (agilex_5_soc_hps2fpga_arready),                                            //  output,   width = 1,                                                                 .arready
		.agilex_5_soc_hps2fpga_rid                                              (agilex_5_soc_hps2fpga_rid),                                                //  output,   width = 4,                                                                 .rid
		.agilex_5_soc_hps2fpga_rdata                                            (agilex_5_soc_hps2fpga_rdata),                                              //  output,  width = 32,                                                                 .rdata
		.agilex_5_soc_hps2fpga_rresp                                            (agilex_5_soc_hps2fpga_rresp),                                              //  output,   width = 2,                                                                 .rresp
		.agilex_5_soc_hps2fpga_rlast                                            (agilex_5_soc_hps2fpga_rlast),                                              //  output,   width = 1,                                                                 .rlast
		.agilex_5_soc_hps2fpga_rvalid                                           (agilex_5_soc_hps2fpga_rvalid),                                             //  output,   width = 1,                                                                 .rvalid
		.agilex_5_soc_hps2fpga_rready                                           (agilex_5_soc_hps2fpga_rready),                                             //   input,   width = 1,                                                                 .rready
		.fpga_only_master_master_address                                        (fpga_only_master_master_address),                                          //   input,  width = 32,                                          fpga_only_master_master.address
		.fpga_only_master_master_waitrequest                                    (fpga_only_master_master_waitrequest),                                      //  output,   width = 1,                                                                 .waitrequest
		.fpga_only_master_master_byteenable                                     (fpga_only_master_master_byteenable),                                       //   input,   width = 4,                                                                 .byteenable
		.fpga_only_master_master_read                                           (fpga_only_master_master_read),                                             //   input,   width = 1,                                                                 .read
		.fpga_only_master_master_readdata                                       (fpga_only_master_master_readdata),                                         //  output,  width = 32,                                                                 .readdata
		.fpga_only_master_master_readdatavalid                                  (fpga_only_master_master_readdatavalid),                                    //  output,   width = 1,                                                                 .readdatavalid
		.fpga_only_master_master_write                                          (fpga_only_master_master_write),                                            //   input,   width = 1,                                                                 .write
		.fpga_only_master_master_writedata                                      (fpga_only_master_master_writedata),                                        //   input,  width = 32,                                                                 .writedata
		.onchip_sram_axi_s1_awid                                                (mm_interconnect_1_onchip_sram_axi_s1_awid),                                //  output,   width = 7,                                               onchip_sram_axi_s1.awid
		.onchip_sram_axi_s1_awaddr                                              (mm_interconnect_1_onchip_sram_axi_s1_awaddr),                              //  output,  width = 15,                                                                 .awaddr
		.onchip_sram_axi_s1_awlen                                               (mm_interconnect_1_onchip_sram_axi_s1_awlen),                               //  output,   width = 8,                                                                 .awlen
		.onchip_sram_axi_s1_awsize                                              (mm_interconnect_1_onchip_sram_axi_s1_awsize),                              //  output,   width = 3,                                                                 .awsize
		.onchip_sram_axi_s1_awburst                                             (mm_interconnect_1_onchip_sram_axi_s1_awburst),                             //  output,   width = 2,                                                                 .awburst
		.onchip_sram_axi_s1_awvalid                                             (mm_interconnect_1_onchip_sram_axi_s1_awvalid),                             //  output,   width = 1,                                                                 .awvalid
		.onchip_sram_axi_s1_awready                                             (mm_interconnect_1_onchip_sram_axi_s1_awready),                             //   input,   width = 1,                                                                 .awready
		.onchip_sram_axi_s1_wdata                                               (mm_interconnect_1_onchip_sram_axi_s1_wdata),                               //  output,  width = 64,                                                                 .wdata
		.onchip_sram_axi_s1_wstrb                                               (mm_interconnect_1_onchip_sram_axi_s1_wstrb),                               //  output,   width = 8,                                                                 .wstrb
		.onchip_sram_axi_s1_wlast                                               (mm_interconnect_1_onchip_sram_axi_s1_wlast),                               //  output,   width = 1,                                                                 .wlast
		.onchip_sram_axi_s1_wvalid                                              (mm_interconnect_1_onchip_sram_axi_s1_wvalid),                              //  output,   width = 1,                                                                 .wvalid
		.onchip_sram_axi_s1_wready                                              (mm_interconnect_1_onchip_sram_axi_s1_wready),                              //   input,   width = 1,                                                                 .wready
		.onchip_sram_axi_s1_bid                                                 (mm_interconnect_1_onchip_sram_axi_s1_bid),                                 //   input,   width = 7,                                                                 .bid
		.onchip_sram_axi_s1_bresp                                               (mm_interconnect_1_onchip_sram_axi_s1_bresp),                               //   input,   width = 2,                                                                 .bresp
		.onchip_sram_axi_s1_bvalid                                              (mm_interconnect_1_onchip_sram_axi_s1_bvalid),                              //   input,   width = 1,                                                                 .bvalid
		.onchip_sram_axi_s1_bready                                              (mm_interconnect_1_onchip_sram_axi_s1_bready),                              //  output,   width = 1,                                                                 .bready
		.onchip_sram_axi_s1_arid                                                (mm_interconnect_1_onchip_sram_axi_s1_arid),                                //  output,   width = 7,                                                                 .arid
		.onchip_sram_axi_s1_araddr                                              (mm_interconnect_1_onchip_sram_axi_s1_araddr),                              //  output,  width = 15,                                                                 .araddr
		.onchip_sram_axi_s1_arlen                                               (mm_interconnect_1_onchip_sram_axi_s1_arlen),                               //  output,   width = 8,                                                                 .arlen
		.onchip_sram_axi_s1_arsize                                              (mm_interconnect_1_onchip_sram_axi_s1_arsize),                              //  output,   width = 3,                                                                 .arsize
		.onchip_sram_axi_s1_arburst                                             (mm_interconnect_1_onchip_sram_axi_s1_arburst),                             //  output,   width = 2,                                                                 .arburst
		.onchip_sram_axi_s1_arvalid                                             (mm_interconnect_1_onchip_sram_axi_s1_arvalid),                             //  output,   width = 1,                                                                 .arvalid
		.onchip_sram_axi_s1_arready                                             (mm_interconnect_1_onchip_sram_axi_s1_arready),                             //   input,   width = 1,                                                                 .arready
		.onchip_sram_axi_s1_rid                                                 (mm_interconnect_1_onchip_sram_axi_s1_rid),                                 //   input,   width = 7,                                                                 .rid
		.onchip_sram_axi_s1_rdata                                               (mm_interconnect_1_onchip_sram_axi_s1_rdata),                               //   input,  width = 64,                                                                 .rdata
		.onchip_sram_axi_s1_rresp                                               (mm_interconnect_1_onchip_sram_axi_s1_rresp),                               //   input,   width = 2,                                                                 .rresp
		.onchip_sram_axi_s1_rlast                                               (mm_interconnect_1_onchip_sram_axi_s1_rlast),                               //   input,   width = 1,                                                                 .rlast
		.onchip_sram_axi_s1_rvalid                                              (mm_interconnect_1_onchip_sram_axi_s1_rvalid),                              //   input,   width = 1,                                                                 .rvalid
		.onchip_sram_axi_s1_rready                                              (mm_interconnect_1_onchip_sram_axi_s1_rready),                              //  output,   width = 1,                                                                 .rready
		.peripheral_sys_0_mm_peripheral_bridge_s0_address                       (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_address),       //  output,  width = 24,                         peripheral_sys_0_mm_peripheral_bridge_s0.address
		.peripheral_sys_0_mm_peripheral_bridge_s0_write                         (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_write),         //  output,   width = 1,                                                                 .write
		.peripheral_sys_0_mm_peripheral_bridge_s0_read                          (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_read),          //  output,   width = 1,                                                                 .read
		.peripheral_sys_0_mm_peripheral_bridge_s0_readdata                      (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_readdata),      //   input,  width = 32,                                                                 .readdata
		.peripheral_sys_0_mm_peripheral_bridge_s0_writedata                     (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_writedata),     //  output,  width = 32,                                                                 .writedata
		.peripheral_sys_0_mm_peripheral_bridge_s0_burstcount                    (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_burstcount),    //  output,   width = 1,                                                                 .burstcount
		.peripheral_sys_0_mm_peripheral_bridge_s0_byteenable                    (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_byteenable),    //  output,   width = 4,                                                                 .byteenable
		.peripheral_sys_0_mm_peripheral_bridge_s0_readdatavalid                 (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_readdatavalid), //   input,   width = 1,                                                                 .readdatavalid
		.peripheral_sys_0_mm_peripheral_bridge_s0_waitrequest                   (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_waitrequest),   //   input,   width = 1,                                                                 .waitrequest
		.peripheral_sys_0_mm_peripheral_bridge_s0_debugaccess                   (mm_interconnect_1_peripheral_sys_0_mm_peripheral_bridge_s0_debugaccess),   //  output,   width = 1,                                                                 .debugaccess
		.onchip_sram_reset1_reset_bridge_in_reset_reset                         (rst_controller_005_reset_out_reset),                                       //   input,   width = 1,                         onchip_sram_reset1_reset_bridge_in_reset.reset
		.peripheral_sys_0_reset_reset_bridge_in_reset_reset                     (rst_controller_004_reset_out_reset),                                       //   input,   width = 1,                     peripheral_sys_0_reset_reset_bridge_in_reset.reset
		.agilex_5_soc_hps2fpga_translator_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                                       //   input,   width = 1, agilex_5_soc_hps2fpga_translator_clk_reset_reset_bridge_in_reset.reset
		.fpga_only_master_master_translator_reset_reset_bridge_in_reset_reset   (rst_controller_006_reset_out_reset),                                       //   input,   width = 1,   fpga_only_master_master_translator_reset_reset_bridge_in_reset.reset
		.onchip_sram_axi_s1_translator_clk_reset_reset_bridge_in_reset_reset    (rst_controller_005_reset_out_reset),                                       //   input,   width = 1,    onchip_sram_axi_s1_translator_clk_reset_reset_bridge_in_reset.reset
		.crosser_002_in_clk_reset_reset_bridge_in_reset_reset                   (rst_controller_006_reset_out_reset),                                       //   input,   width = 1,                   crosser_002_in_clk_reset_reset_bridge_in_reset.reset
		.agilex_5_soc_h2f_user1_clk_clk                                         (agilex_5_soc_h2f_user1_clk_clk),                                           //   input,   width = 1,                                       agilex_5_soc_h2f_user1_clk.clk
		.agilex_5_soc_h2f_user0_clk_clk                                         (agilex_5_soc_h2f_user0_clk_clk)                                            //   input,   width = 1,                                       agilex_5_soc_h2f_user0_clk.clk
	);

	ghrd_hps_system_altera_mm_interconnect_1920_fivhe3y mm_interconnect_2 (
		.agilex_5_soc_lwhps2fpga_awid                                             (agilex_5_soc_lwhps2fpga_awid),                                   //   input,   width = 4,                                            agilex_5_soc_lwhps2fpga.awid
		.agilex_5_soc_lwhps2fpga_awaddr                                           (agilex_5_soc_lwhps2fpga_awaddr),                                 //   input,  width = 29,                                                                   .awaddr
		.agilex_5_soc_lwhps2fpga_awlen                                            (agilex_5_soc_lwhps2fpga_awlen),                                  //   input,   width = 8,                                                                   .awlen
		.agilex_5_soc_lwhps2fpga_awsize                                           (agilex_5_soc_lwhps2fpga_awsize),                                 //   input,   width = 3,                                                                   .awsize
		.agilex_5_soc_lwhps2fpga_awburst                                          (agilex_5_soc_lwhps2fpga_awburst),                                //   input,   width = 2,                                                                   .awburst
		.agilex_5_soc_lwhps2fpga_awlock                                           (agilex_5_soc_lwhps2fpga_awlock),                                 //   input,   width = 1,                                                                   .awlock
		.agilex_5_soc_lwhps2fpga_awcache                                          (agilex_5_soc_lwhps2fpga_awcache),                                //   input,   width = 4,                                                                   .awcache
		.agilex_5_soc_lwhps2fpga_awprot                                           (agilex_5_soc_lwhps2fpga_awprot),                                 //   input,   width = 3,                                                                   .awprot
		.agilex_5_soc_lwhps2fpga_awvalid                                          (agilex_5_soc_lwhps2fpga_awvalid),                                //   input,   width = 1,                                                                   .awvalid
		.agilex_5_soc_lwhps2fpga_awready                                          (agilex_5_soc_lwhps2fpga_awready),                                //  output,   width = 1,                                                                   .awready
		.agilex_5_soc_lwhps2fpga_wdata                                            (agilex_5_soc_lwhps2fpga_wdata),                                  //   input,  width = 32,                                                                   .wdata
		.agilex_5_soc_lwhps2fpga_wstrb                                            (agilex_5_soc_lwhps2fpga_wstrb),                                  //   input,   width = 4,                                                                   .wstrb
		.agilex_5_soc_lwhps2fpga_wlast                                            (agilex_5_soc_lwhps2fpga_wlast),                                  //   input,   width = 1,                                                                   .wlast
		.agilex_5_soc_lwhps2fpga_wvalid                                           (agilex_5_soc_lwhps2fpga_wvalid),                                 //   input,   width = 1,                                                                   .wvalid
		.agilex_5_soc_lwhps2fpga_wready                                           (agilex_5_soc_lwhps2fpga_wready),                                 //  output,   width = 1,                                                                   .wready
		.agilex_5_soc_lwhps2fpga_bid                                              (agilex_5_soc_lwhps2fpga_bid),                                    //  output,   width = 4,                                                                   .bid
		.agilex_5_soc_lwhps2fpga_bresp                                            (agilex_5_soc_lwhps2fpga_bresp),                                  //  output,   width = 2,                                                                   .bresp
		.agilex_5_soc_lwhps2fpga_bvalid                                           (agilex_5_soc_lwhps2fpga_bvalid),                                 //  output,   width = 1,                                                                   .bvalid
		.agilex_5_soc_lwhps2fpga_bready                                           (agilex_5_soc_lwhps2fpga_bready),                                 //   input,   width = 1,                                                                   .bready
		.agilex_5_soc_lwhps2fpga_arid                                             (agilex_5_soc_lwhps2fpga_arid),                                   //   input,   width = 4,                                                                   .arid
		.agilex_5_soc_lwhps2fpga_araddr                                           (agilex_5_soc_lwhps2fpga_araddr),                                 //   input,  width = 29,                                                                   .araddr
		.agilex_5_soc_lwhps2fpga_arlen                                            (agilex_5_soc_lwhps2fpga_arlen),                                  //   input,   width = 8,                                                                   .arlen
		.agilex_5_soc_lwhps2fpga_arsize                                           (agilex_5_soc_lwhps2fpga_arsize),                                 //   input,   width = 3,                                                                   .arsize
		.agilex_5_soc_lwhps2fpga_arburst                                          (agilex_5_soc_lwhps2fpga_arburst),                                //   input,   width = 2,                                                                   .arburst
		.agilex_5_soc_lwhps2fpga_arlock                                           (agilex_5_soc_lwhps2fpga_arlock),                                 //   input,   width = 1,                                                                   .arlock
		.agilex_5_soc_lwhps2fpga_arcache                                          (agilex_5_soc_lwhps2fpga_arcache),                                //   input,   width = 4,                                                                   .arcache
		.agilex_5_soc_lwhps2fpga_arprot                                           (agilex_5_soc_lwhps2fpga_arprot),                                 //   input,   width = 3,                                                                   .arprot
		.agilex_5_soc_lwhps2fpga_arvalid                                          (agilex_5_soc_lwhps2fpga_arvalid),                                //   input,   width = 1,                                                                   .arvalid
		.agilex_5_soc_lwhps2fpga_arready                                          (agilex_5_soc_lwhps2fpga_arready),                                //  output,   width = 1,                                                                   .arready
		.agilex_5_soc_lwhps2fpga_rid                                              (agilex_5_soc_lwhps2fpga_rid),                                    //  output,   width = 4,                                                                   .rid
		.agilex_5_soc_lwhps2fpga_rdata                                            (agilex_5_soc_lwhps2fpga_rdata),                                  //  output,  width = 32,                                                                   .rdata
		.agilex_5_soc_lwhps2fpga_rresp                                            (agilex_5_soc_lwhps2fpga_rresp),                                  //  output,   width = 2,                                                                   .rresp
		.agilex_5_soc_lwhps2fpga_rlast                                            (agilex_5_soc_lwhps2fpga_rlast),                                  //  output,   width = 1,                                                                   .rlast
		.agilex_5_soc_lwhps2fpga_rvalid                                           (agilex_5_soc_lwhps2fpga_rvalid),                                 //  output,   width = 1,                                                                   .rvalid
		.agilex_5_soc_lwhps2fpga_rready                                           (agilex_5_soc_lwhps2fpga_rready),                                 //   input,   width = 1,                                                                   .rready
		.video_sys_0_mm_video_bridge_s0_address                                   (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_address),       //  output,  width = 24,                                     video_sys_0_mm_video_bridge_s0.address
		.video_sys_0_mm_video_bridge_s0_write                                     (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_write),         //  output,   width = 1,                                                                   .write
		.video_sys_0_mm_video_bridge_s0_read                                      (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_read),          //  output,   width = 1,                                                                   .read
		.video_sys_0_mm_video_bridge_s0_readdata                                  (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_readdata),      //   input,  width = 32,                                                                   .readdata
		.video_sys_0_mm_video_bridge_s0_writedata                                 (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_writedata),     //  output,  width = 32,                                                                   .writedata
		.video_sys_0_mm_video_bridge_s0_burstcount                                (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_burstcount),    //  output,   width = 1,                                                                   .burstcount
		.video_sys_0_mm_video_bridge_s0_byteenable                                (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_byteenable),    //  output,   width = 4,                                                                   .byteenable
		.video_sys_0_mm_video_bridge_s0_readdatavalid                             (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_readdatavalid), //   input,   width = 1,                                                                   .readdatavalid
		.video_sys_0_mm_video_bridge_s0_waitrequest                               (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_waitrequest),   //   input,   width = 1,                                                                   .waitrequest
		.video_sys_0_mm_video_bridge_s0_debugaccess                               (mm_interconnect_2_video_sys_0_mm_video_bridge_s0_debugaccess),   //  output,   width = 1,                                                                   .debugaccess
		.emif_bank3a_s0_axil_awaddr                                               (mm_interconnect_2_emif_bank3a_s0_axil_awaddr),                   //  output,  width = 27,                                                emif_bank3a_s0_axil.awaddr
		.emif_bank3a_s0_axil_awprot                                               (mm_interconnect_2_emif_bank3a_s0_axil_awprot),                   //  output,   width = 3,                                                                   .awprot
		.emif_bank3a_s0_axil_awvalid                                              (mm_interconnect_2_emif_bank3a_s0_axil_awvalid),                  //  output,   width = 1,                                                                   .awvalid
		.emif_bank3a_s0_axil_awready                                              (mm_interconnect_2_emif_bank3a_s0_axil_awready),                  //   input,   width = 1,                                                                   .awready
		.emif_bank3a_s0_axil_wdata                                                (mm_interconnect_2_emif_bank3a_s0_axil_wdata),                    //  output,  width = 32,                                                                   .wdata
		.emif_bank3a_s0_axil_wstrb                                                (mm_interconnect_2_emif_bank3a_s0_axil_wstrb),                    //  output,   width = 4,                                                                   .wstrb
		.emif_bank3a_s0_axil_wvalid                                               (mm_interconnect_2_emif_bank3a_s0_axil_wvalid),                   //  output,   width = 1,                                                                   .wvalid
		.emif_bank3a_s0_axil_wready                                               (mm_interconnect_2_emif_bank3a_s0_axil_wready),                   //   input,   width = 1,                                                                   .wready
		.emif_bank3a_s0_axil_bresp                                                (mm_interconnect_2_emif_bank3a_s0_axil_bresp),                    //   input,   width = 2,                                                                   .bresp
		.emif_bank3a_s0_axil_bvalid                                               (mm_interconnect_2_emif_bank3a_s0_axil_bvalid),                   //   input,   width = 1,                                                                   .bvalid
		.emif_bank3a_s0_axil_bready                                               (mm_interconnect_2_emif_bank3a_s0_axil_bready),                   //  output,   width = 1,                                                                   .bready
		.emif_bank3a_s0_axil_araddr                                               (mm_interconnect_2_emif_bank3a_s0_axil_araddr),                   //  output,  width = 27,                                                                   .araddr
		.emif_bank3a_s0_axil_arprot                                               (mm_interconnect_2_emif_bank3a_s0_axil_arprot),                   //  output,   width = 3,                                                                   .arprot
		.emif_bank3a_s0_axil_arvalid                                              (mm_interconnect_2_emif_bank3a_s0_axil_arvalid),                  //  output,   width = 1,                                                                   .arvalid
		.emif_bank3a_s0_axil_arready                                              (mm_interconnect_2_emif_bank3a_s0_axil_arready),                  //   input,   width = 1,                                                                   .arready
		.emif_bank3a_s0_axil_rdata                                                (mm_interconnect_2_emif_bank3a_s0_axil_rdata),                    //   input,  width = 32,                                                                   .rdata
		.emif_bank3a_s0_axil_rresp                                                (mm_interconnect_2_emif_bank3a_s0_axil_rresp),                    //   input,   width = 2,                                                                   .rresp
		.emif_bank3a_s0_axil_rvalid                                               (mm_interconnect_2_emif_bank3a_s0_axil_rvalid),                   //   input,   width = 1,                                                                   .rvalid
		.emif_bank3a_s0_axil_rready                                               (mm_interconnect_2_emif_bank3a_s0_axil_rready),                   //  output,   width = 1,                                                                   .rready
		.video_sys_0_reset_reset_bridge_in_reset_reset                            (rst_controller_004_reset_out_reset),                             //   input,   width = 1,                            video_sys_0_reset_reset_bridge_in_reset.reset
		.agilex_5_soc_lwhps2fpga_translator_clk_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),                             //   input,   width = 1, agilex_5_soc_lwhps2fpga_translator_clk_reset_reset_bridge_in_reset.reset
		.emif_bank3a_s0_axil_agent_reset_sink_reset_bridge_in_reset_reset         (rst_controller_007_reset_out_reset),                             //   input,   width = 1,         emif_bank3a_s0_axil_agent_reset_sink_reset_bridge_in_reset.reset
		.agilex_5_soc_h2f_user1_clk_clk                                           (agilex_5_soc_h2f_user1_clk_clk)                                  //   input,   width = 1,                                         agilex_5_soc_h2f_user1_clk.clk
	);

	ghrd_hps_system_altera_mm_interconnect_1920_xvazuei mm_interconnect_3 (
		.bank3a_emif_master_master_address                                      (bank3a_emif_master_master_address),             //   input,   width = 32,                                        bank3a_emif_master_master.address
		.bank3a_emif_master_master_waitrequest                                  (bank3a_emif_master_master_waitrequest),         //  output,    width = 1,                                                                 .waitrequest
		.bank3a_emif_master_master_byteenable                                   (bank3a_emif_master_master_byteenable),          //   input,    width = 4,                                                                 .byteenable
		.bank3a_emif_master_master_read                                         (bank3a_emif_master_master_read),                //   input,    width = 1,                                                                 .read
		.bank3a_emif_master_master_readdata                                     (bank3a_emif_master_master_readdata),            //  output,   width = 32,                                                                 .readdata
		.bank3a_emif_master_master_readdatavalid                                (bank3a_emif_master_master_readdatavalid),       //  output,    width = 1,                                                                 .readdatavalid
		.bank3a_emif_master_master_write                                        (bank3a_emif_master_master_write),               //   input,    width = 1,                                                                 .write
		.bank3a_emif_master_master_writedata                                    (bank3a_emif_master_master_writedata),           //   input,   width = 32,                                                                 .writedata
		.emif_bank3a_s0_axi4_awid                                               (mm_interconnect_3_emif_bank3a_s0_axi4_awid),    //  output,    width = 7,                                              emif_bank3a_s0_axi4.awid
		.emif_bank3a_s0_axi4_awaddr                                             (mm_interconnect_3_emif_bank3a_s0_axi4_awaddr),  //  output,   width = 32,                                                                 .awaddr
		.emif_bank3a_s0_axi4_awlen                                              (mm_interconnect_3_emif_bank3a_s0_axi4_awlen),   //  output,    width = 8,                                                                 .awlen
		.emif_bank3a_s0_axi4_awsize                                             (mm_interconnect_3_emif_bank3a_s0_axi4_awsize),  //  output,    width = 3,                                                                 .awsize
		.emif_bank3a_s0_axi4_awburst                                            (mm_interconnect_3_emif_bank3a_s0_axi4_awburst), //  output,    width = 2,                                                                 .awburst
		.emif_bank3a_s0_axi4_awlock                                             (mm_interconnect_3_emif_bank3a_s0_axi4_awlock),  //  output,    width = 1,                                                                 .awlock
		.emif_bank3a_s0_axi4_awprot                                             (mm_interconnect_3_emif_bank3a_s0_axi4_awprot),  //  output,    width = 3,                                                                 .awprot
		.emif_bank3a_s0_axi4_awuser                                             (mm_interconnect_3_emif_bank3a_s0_axi4_awuser),  //  output,   width = 14,                                                                 .awuser
		.emif_bank3a_s0_axi4_awqos                                              (mm_interconnect_3_emif_bank3a_s0_axi4_awqos),   //  output,    width = 4,                                                                 .awqos
		.emif_bank3a_s0_axi4_awvalid                                            (mm_interconnect_3_emif_bank3a_s0_axi4_awvalid), //  output,    width = 1,                                                                 .awvalid
		.emif_bank3a_s0_axi4_awready                                            (mm_interconnect_3_emif_bank3a_s0_axi4_awready), //   input,    width = 1,                                                                 .awready
		.emif_bank3a_s0_axi4_wdata                                              (mm_interconnect_3_emif_bank3a_s0_axi4_wdata),   //  output,  width = 256,                                                                 .wdata
		.emif_bank3a_s0_axi4_wstrb                                              (mm_interconnect_3_emif_bank3a_s0_axi4_wstrb),   //  output,   width = 32,                                                                 .wstrb
		.emif_bank3a_s0_axi4_wlast                                              (mm_interconnect_3_emif_bank3a_s0_axi4_wlast),   //  output,    width = 1,                                                                 .wlast
		.emif_bank3a_s0_axi4_wvalid                                             (mm_interconnect_3_emif_bank3a_s0_axi4_wvalid),  //  output,    width = 1,                                                                 .wvalid
		.emif_bank3a_s0_axi4_wuser                                              (mm_interconnect_3_emif_bank3a_s0_axi4_wuser),   //  output,   width = 64,                                                                 .wuser
		.emif_bank3a_s0_axi4_wready                                             (mm_interconnect_3_emif_bank3a_s0_axi4_wready),  //   input,    width = 1,                                                                 .wready
		.emif_bank3a_s0_axi4_bid                                                (mm_interconnect_3_emif_bank3a_s0_axi4_bid),     //   input,    width = 7,                                                                 .bid
		.emif_bank3a_s0_axi4_bresp                                              (mm_interconnect_3_emif_bank3a_s0_axi4_bresp),   //   input,    width = 2,                                                                 .bresp
		.emif_bank3a_s0_axi4_bvalid                                             (mm_interconnect_3_emif_bank3a_s0_axi4_bvalid),  //   input,    width = 1,                                                                 .bvalid
		.emif_bank3a_s0_axi4_bready                                             (mm_interconnect_3_emif_bank3a_s0_axi4_bready),  //  output,    width = 1,                                                                 .bready
		.emif_bank3a_s0_axi4_arid                                               (mm_interconnect_3_emif_bank3a_s0_axi4_arid),    //  output,    width = 7,                                                                 .arid
		.emif_bank3a_s0_axi4_araddr                                             (mm_interconnect_3_emif_bank3a_s0_axi4_araddr),  //  output,   width = 32,                                                                 .araddr
		.emif_bank3a_s0_axi4_arlen                                              (mm_interconnect_3_emif_bank3a_s0_axi4_arlen),   //  output,    width = 8,                                                                 .arlen
		.emif_bank3a_s0_axi4_arsize                                             (mm_interconnect_3_emif_bank3a_s0_axi4_arsize),  //  output,    width = 3,                                                                 .arsize
		.emif_bank3a_s0_axi4_arburst                                            (mm_interconnect_3_emif_bank3a_s0_axi4_arburst), //  output,    width = 2,                                                                 .arburst
		.emif_bank3a_s0_axi4_arlock                                             (mm_interconnect_3_emif_bank3a_s0_axi4_arlock),  //  output,    width = 1,                                                                 .arlock
		.emif_bank3a_s0_axi4_arprot                                             (mm_interconnect_3_emif_bank3a_s0_axi4_arprot),  //  output,    width = 3,                                                                 .arprot
		.emif_bank3a_s0_axi4_aruser                                             (mm_interconnect_3_emif_bank3a_s0_axi4_aruser),  //  output,   width = 14,                                                                 .aruser
		.emif_bank3a_s0_axi4_arqos                                              (mm_interconnect_3_emif_bank3a_s0_axi4_arqos),   //  output,    width = 4,                                                                 .arqos
		.emif_bank3a_s0_axi4_arvalid                                            (mm_interconnect_3_emif_bank3a_s0_axi4_arvalid), //  output,    width = 1,                                                                 .arvalid
		.emif_bank3a_s0_axi4_arready                                            (mm_interconnect_3_emif_bank3a_s0_axi4_arready), //   input,    width = 1,                                                                 .arready
		.emif_bank3a_s0_axi4_rid                                                (mm_interconnect_3_emif_bank3a_s0_axi4_rid),     //   input,    width = 7,                                                                 .rid
		.emif_bank3a_s0_axi4_rdata                                              (mm_interconnect_3_emif_bank3a_s0_axi4_rdata),   //   input,  width = 256,                                                                 .rdata
		.emif_bank3a_s0_axi4_rresp                                              (mm_interconnect_3_emif_bank3a_s0_axi4_rresp),   //   input,    width = 2,                                                                 .rresp
		.emif_bank3a_s0_axi4_rlast                                              (mm_interconnect_3_emif_bank3a_s0_axi4_rlast),   //   input,    width = 1,                                                                 .rlast
		.emif_bank3a_s0_axi4_rvalid                                             (mm_interconnect_3_emif_bank3a_s0_axi4_rvalid),  //   input,    width = 1,                                                                 .rvalid
		.emif_bank3a_s0_axi4_rready                                             (mm_interconnect_3_emif_bank3a_s0_axi4_rready),  //  output,    width = 1,                                                                 .rready
		.emif_bank3a_s0_axi4_ruser                                              (mm_interconnect_3_emif_bank3a_s0_axi4_ruser),   //   input,   width = 64,                                                                 .ruser
		.bank3a_emif_master_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),            //   input,    width = 1, bank3a_emif_master_master_translator_reset_reset_bridge_in_reset.reset
		.emif_bank3a_s0_axi4_translator_clk_reset_reset_bridge_in_reset_reset   (rst_controller_008_reset_out_reset),            //   input,    width = 1,   emif_bank3a_s0_axi4_translator_clk_reset_reset_bridge_in_reset.reset
		.agilex_5_soc_h2f_user1_clk_clk                                         (agilex_5_soc_h2f_user1_clk_clk)                 //   input,    width = 1,                                       agilex_5_soc_h2f_user1_clk.clk
	);

	ghrd_hps_system_altera_irq_mapper_2000_3dsv57y irq_mapper (
		.clk           (),                                    //   input,   width = 1,       clk.clk
		.reset         (),                                    //   input,   width = 1, clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),            //   input,   width = 1, receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),            //   input,   width = 1, receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),            //   input,   width = 1, receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),            //   input,   width = 1, receiver3.irq
		.sender_irq    (agilex_5_soc_fpga2hps_interrupt_irq)  //  output,  width = 63,    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~agilex_5_soc_h2f_cold_reset_reset), //   input,  width = 1, reset_in0.reset
		.reset_in1      (~agilex_5_soc_h2f_reset_reset),      //   input,  width = 1, reset_in1.reset
		.clk            (),                                   //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~agilex_5_soc_h2f_cold_reset_reset), //   input,  width = 1, reset_in0.reset
		.reset_in1      (~agilex_5_soc_h2f_reset_reset),      //   input,  width = 1, reset_in1.reset
		.clk            (agilex_5_soc_h2f_user1_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (fpga_only_master_master_reset_reset), //   input,  width = 1, reset_in0.reset
		.reset_in1      (reset_in_out_reset_reset),            //   input,  width = 1, reset_in1.reset
		.clk            (),                                    //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (reset_in_out_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (agilex_5_soc_h2f_user0_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (reset_in_out_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (agilex_5_soc_h2f_user1_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (reset_in_out_reset_reset),           //   input,  width = 1, reset_in0.reset
		.clk            (agilex_5_soc_h2f_user0_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (fpga_only_master_master_reset_reset), //   input,  width = 1, reset_in0.reset
		.reset_in1      (reset_in_out_reset_reset),            //   input,  width = 1, reset_in1.reset
		.clk            (agilex_5_soc_h2f_user1_clk_clk),      //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                    // (terminated),                       
		.reset_req_in0  (1'b0),                                // (terminated),                       
		.reset_req_in1  (1'b0),                                // (terminated),                       
		.reset_in2      (1'b0),                                // (terminated),                       
		.reset_req_in2  (1'b0),                                // (terminated),                       
		.reset_in3      (1'b0),                                // (terminated),                       
		.reset_req_in3  (1'b0),                                // (terminated),                       
		.reset_in4      (1'b0),                                // (terminated),                       
		.reset_req_in4  (1'b0),                                // (terminated),                       
		.reset_in5      (1'b0),                                // (terminated),                       
		.reset_req_in5  (1'b0),                                // (terminated),                       
		.reset_in6      (1'b0),                                // (terminated),                       
		.reset_req_in6  (1'b0),                                // (terminated),                       
		.reset_in7      (1'b0),                                // (terminated),                       
		.reset_req_in7  (1'b0),                                // (terminated),                       
		.reset_in8      (1'b0),                                // (terminated),                       
		.reset_req_in8  (1'b0),                                // (terminated),                       
		.reset_in9      (1'b0),                                // (terminated),                       
		.reset_req_in9  (1'b0),                                // (terminated),                       
		.reset_in10     (1'b0),                                // (terminated),                       
		.reset_req_in10 (1'b0),                                // (terminated),                       
		.reset_in11     (1'b0),                                // (terminated),                       
		.reset_req_in11 (1'b0),                                // (terminated),                       
		.reset_in12     (1'b0),                                // (terminated),                       
		.reset_req_in12 (1'b0),                                // (terminated),                       
		.reset_in13     (1'b0),                                // (terminated),                       
		.reset_req_in13 (1'b0),                                // (terminated),                       
		.reset_in14     (1'b0),                                // (terminated),                       
		.reset_req_in14 (1'b0),                                // (terminated),                       
		.reset_in15     (1'b0),                                // (terminated),                       
		.reset_req_in15 (1'b0)                                 // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~agilex_5_soc_h2f_cold_reset_reset), //   input,  width = 1, reset_in0.reset
		.reset_in1      (~agilex_5_soc_h2f_reset_reset),      //   input,  width = 1, reset_in1.reset
		.clk            (agilex_5_soc_h2f_user1_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~emif_bank3a_usr_rst_n_0_reset),     //   input,  width = 1, reset_in0.reset
		.clk            (agilex_5_soc_h2f_user1_clk_clk),     //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
