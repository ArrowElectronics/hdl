
module adrv9001_gpio_in (
	ck,
	dout,
	pad_in);	

	input		ck;
	output	[1:0]	dout;
	input	[0:0]	pad_in;
endmodule
