
module input_buf (
	dout,
	pad_in,
	pad_in_b);	

	output	[0:0]	dout;
	input	[0:0]	pad_in;
	input	[0:0]	pad_in_b;
endmodule
