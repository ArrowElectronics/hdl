
module adrv9002_gpio_in (
	dout,
	pad_in,
	ck);	

	output	[1:0]	dout;
	input	[0:0]	pad_in;
	input		ck;
endmodule
