
module adrv9002_gpio_out (
	din,
	pad_out,
	ck);	

	input	[1:0]	din;
	output	[0:0]	pad_out;
	input		ck;
endmodule
